-----------------------------------------------------------------
-- Created By: Richard Cho
-- Create Date: 3/17/2022
-----------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity SCORE_CALC is
    
    port (
        clk : in std_logic; -- system clock
        rst : in std_logic; -- system reset
		temp : in std_logic_vector (8 downto 0); -- celcius
		eda : in std_logic_vector (6 downto 0); --micro siemens
		hr : in std_logic_vector (10 downto 0); -- bpm
		stress_score : out std_logic_vector (47 downto 0); -- output
		not_stress_score : out std_logic_vector (48 downto 0); -- output
		status : out std_logic_vector (1 downto 0)); -- output
		
end SCORE_CALC;

architecture behavioral of SCORE_CALC is

	signal P_TEMP_S : unsigned(11 downto 0);
	signal P_TEMP_NS : unsigned(11 downto 0);
	
	signal P_EDA_S : unsigned(11 downto 0);
	signal P_EDA_NS : unsigned(11 downto 0);
	
	signal P_HR_S : unsigned(11 downto 0);
	signal P_HR_NS : unsigned(11 downto 0);
	
	signal stress_score_temp : unsigned(47 downto 0);
	signal not_stress_score_temp : unsigned(48 downto 0);
	
	-- constants
	constant P_STRESS : unsigned(11 downto 0) := "011111010000";
	constant P_NOT_STRESS : unsigned(12 downto 0) := "1111101000000";
	
begin
	process(temp, eda, hr) -- stress score
	begin
		case temp is
			when "011111110" => P_TEMP_S <= "001101100000";
			when "011111111" => P_TEMP_S <= "100100101111";
			when "100000000" => P_TEMP_S <= "001110100010";
			when "100000001" => P_TEMP_S <= "010000010010";
			when "100000010" => P_TEMP_S <= "001001111100";
			when "100000011" => P_TEMP_S <= "000100001010";
			when "100000100" => P_TEMP_S <= "000010111001";
			when "100000101" => P_TEMP_S <= "000010100101";
			when "100000110" => P_TEMP_S <= "000010011100";
			when "100000111" => P_TEMP_S <= "000010100001";
			when "100001000" => P_TEMP_S <= "000010010110";
			when "100001001" => P_TEMP_S <= "000010001011";
			when "100001010" => P_TEMP_S <= "000010100000";
			when "100001011" => P_TEMP_S <= "000111100100";
			when "100001100" => P_TEMP_S <= "001000001110";
			when "100001101" => P_TEMP_S <= "001001001001";
			when "100001110" => P_TEMP_S <= "000011111011";
			when "100001111" => P_TEMP_S <= "000100111110";
			when "100010000" => P_TEMP_S <= "000001101100";
			when "100010001" => P_TEMP_S <= "000001110110";
			when "100010010" => P_TEMP_S <= "000010010111";
			when "100010011" => P_TEMP_S <= "000011111001";
			when "100010100" => P_TEMP_S <= "000000000010";
			when others => P_TEMP_S      <= "000000000001";
		end case;
		
		case eda is
			when "0110111" => P_EDA_S <= "001001000011";
			when "0111000" => P_EDA_S <= "000101010010";
			when "0111001" => P_EDA_S <= "000000101111";
			when "0111010" => P_EDA_S <= "000010111111";
			when "0111011" => P_EDA_S <= "000101010011";
			when "0111100" => P_EDA_S <= "001000001111";
			when "0111101" => P_EDA_S <= "000101110001";
			when "0111110" => P_EDA_S <= "001011010011";
			when "0111111" => P_EDA_S <= "001100110110";
			when "1000000" => P_EDA_S <= "000111111110";
			when "1000001" => P_EDA_S <= "001010111101";
			when "1000010" => P_EDA_S <= "001001110101";
			when "1000011" => P_EDA_S <= "001000010001";
			when "1000100" => P_EDA_S <= "000111110101";
			when "1000101" => P_EDA_S <= "000011110010";
			when "1000110" => P_EDA_S <= "000101010101";
			when "1000111" => P_EDA_S <= "000011001110";
			when "1001000" => P_EDA_S <= "000011011010";
			when "1001001" => P_EDA_S <= "000010101000";
			when "1001010" => P_EDA_S <= "000011101000";
			when "1001011" => P_EDA_S <= "000011111001";
			when "1001100" => P_EDA_S <= "001010001000";
			when "1001101" => P_EDA_S <= "000011001100";
			when "1001110" => P_EDA_S <= "000000001010";
			when "1001111" | "1010000" => P_EDA_S <= "000000001000";
			when "1010001" => P_EDA_S <= "000000010110";
			when "1010010" => P_EDA_S <= "000000100011";
			when "1010011" | "1011100" => P_EDA_S <= "000000011010";
			when "1010100" | "1011001" => P_EDA_S <= "000000011100";
			when "1010101" => P_EDA_S <= "000000111110";
			when "1010110" => P_EDA_S <= "000001001011";
			when "1010111" => P_EDA_S <= "000001000000";
			when "1011000" | "1011011" => P_EDA_S <= "000000111010";
			when "1011010" => P_EDA_S <= "000000100110";
			when "1011101" => P_EDA_S <= "000000010000";
			when "1011110" => P_EDA_S <= "000000011000";
			when "1011111" => P_EDA_S <= "000001000011";
			when "1100000" => P_EDA_S <= "000000100001";
			when others    => P_EDA_S <= "000000000001";
		end case;

		case hr is
			when "00110010011" => P_HR_S <= "000000001011";
			when "00110010111" => P_HR_S <= "000000001011";
			when "00110011000" => P_HR_S <= "000000001011";
			when "00110011001" => P_HR_S <= "000000001011";
			when "00110110011" => P_HR_S <= "000000010110";
			when "00110110110" => P_HR_S <= "000000001011";
			when "00110111100" => P_HR_S <= "000000010110";
			when "00110111110" => P_HR_S <= "000000001011";
			when "00111000000" => P_HR_S <= "000000001011";
			when "00111000010" => P_HR_S <= "000000001011";
			when "00111000011" => P_HR_S <= "000000001011";
			when "00111000111" => P_HR_S <= "000000010110";
			when "00111001001" => P_HR_S <= "000000010110";
			when "00111001100" => P_HR_S <= "000000001011";
			when "00111001101" => P_HR_S <= "000000001011";
			when "00111001111" => P_HR_S <= "000000001011";
			when "00111010010" => P_HR_S <= "000000001011";
			when "00111010101" => P_HR_S <= "000000001011";
			when "00111010111" => P_HR_S <= "000000001011";
			when "00111011000" => P_HR_S <= "000000001011";
			when "00111011001" => P_HR_S <= "000000001011";
			when "00111011100" => P_HR_S <= "000000100001";
			when "00111011101" => P_HR_S <= "000000100001";
			when "00111100001" => P_HR_S <= "000000100001";
			when "00111100011" => P_HR_S <= "000000001011";
			when "00111100110" => P_HR_S <= "000000001011";
			when "00111101011" => P_HR_S <= "000000001011";
			when "00111101111" => P_HR_S <= "000000010110";
			when "00111110000" => P_HR_S <= "000000001011";
			when "00111110010" => P_HR_S <= "000000001011";
			when "00111110100" => P_HR_S <= "000000001011";
			when "00111110101" => P_HR_S <= "000000010110";
			when "00111110110" => P_HR_S <= "000000010110";
			when "00111111000" => P_HR_S <= "000000001011";
			when "00111111001" => P_HR_S <= "000000010110";
			when "00111111100" => P_HR_S <= "000000010110";
			when "01000000100" => P_HR_S <= "000000010110";
			when "01000000101" => P_HR_S <= "000000001011";
			when "01000000110" => P_HR_S <= "000000010110";
			when "01000000111" => P_HR_S <= "000000010110";
			when "01000001001" => P_HR_S <= "000000001011";
			when "01000001010" => P_HR_S <= "000000001011";
			when "01000001011" => P_HR_S <= "000000001011";
			when "01000001101" => P_HR_S <= "000000001011";
			when "01000001111" => P_HR_S <= "000000101011";
			when "01000010001" => P_HR_S <= "000000101011";
			when "01000010010" => P_HR_S <= "000000010110";
			when "01000010100" => P_HR_S <= "000000110110";
			when "01000010101" => P_HR_S <= "000000001011";
			when "01000010110" => P_HR_S <= "000000010110";
			when "01000010111" => P_HR_S <= "000000001011";
			when "01000011010" => P_HR_S <= "000000101011";
			when "01000011011" => P_HR_S <= "000000100001";
			when "01000011100" => P_HR_S <= "000000001011";
			when "01000011101" => P_HR_S <= "000000001011";
			when "01000100001" => P_HR_S <= "000000100001";
			when "01000100011" => P_HR_S <= "000000001011";
			when "01000100100" => P_HR_S <= "000000001011";
			when "01000100111" => P_HR_S <= "000000001011";
			when "01000101000" => P_HR_S <= "000000010110";
			when "01000101001" => P_HR_S <= "000000001011";
			when "01000101010" => P_HR_S <= "000000101011";
			when "01000101011" => P_HR_S <= "000000110110";
			when "01000101100" => P_HR_S <= "000000010110";
			when "01000101101" => P_HR_S <= "000000010110";
			when "01000101110" => P_HR_S <= "000000001011";
			when "01000101111" => P_HR_S <= "000000100001";
			when "01000110011" => P_HR_S <= "000000100001";
			when "01000110110" => P_HR_S <= "000000010110";
			when "01000110111" => P_HR_S <= "000000001011";
			when "01000111000" => P_HR_S <= "000000010110";
			when "01000111001" => P_HR_S <= "000001001100";
			when "01000111010" => P_HR_S <= "000000010110";
			when "01000111011" => P_HR_S <= "000000001011";
			when "01000111100" => P_HR_S <= "000000001011";
			when "01000111101" => P_HR_S <= "000000100001";
			when "01000111110" => P_HR_S <= "000000100001";
			when "01000111111" => P_HR_S <= "000000010110";
			when "01001000000" => P_HR_S <= "000000001011";
			when "01001000010" => P_HR_S <= "000000101011";
			when "01001000011" => P_HR_S <= "000000001011";
			when "01001000100" => P_HR_S <= "000000101011";
			when "01001000101" => P_HR_S <= "000000010110";
			when "01001000110" => P_HR_S <= "000000001011";
			when "01001000111" => P_HR_S <= "000000100001";
			when "01001001001" => P_HR_S <= "000000100001";
			when "01001001010" => P_HR_S <= "000000010110";
			when "01001001011" => P_HR_S <= "000000100001";
			when "01001001100" => P_HR_S <= "000000001011";
			when "01001001101" => P_HR_S <= "000000110110";
			when "01001010001" => P_HR_S <= "000000010110";
			when "01001010010" => P_HR_S <= "000000001011";
			when "01001010011" => P_HR_S <= "000000001011";
			when "01001010100" => P_HR_S <= "000000101011";
			when "01001010101" => P_HR_S <= "000000001011";
			when "01001010110" => P_HR_S <= "000000100001";
			when "01001010111" => P_HR_S <= "000000001011";
			when "01001011001" => P_HR_S <= "000000001011";
			when "01001011010" => P_HR_S <= "000000100001";
			when "01001011011" => P_HR_S <= "000000010110";
			when "01001011101" => P_HR_S <= "000000101011";
			when "01001011110" => P_HR_S <= "000000101011";
			when "01001100001" => P_HR_S <= "000000010110";
			when "01001100010" => P_HR_S <= "000000100001";
			when "01001100011" => P_HR_S <= "000000010110";
			when "01001100100" => P_HR_S <= "000000010110";
			when "01001100101" => P_HR_S <= "000000010110";
			when "01001100110" => P_HR_S <= "000000100001";
			when "01001100111" => P_HR_S <= "000000010110";
			when "01001101001" => P_HR_S <= "000000001011";
			when "01001101010" => P_HR_S <= "000000001011";
			when "01001101011" => P_HR_S <= "000000110110";
			when "01001101100" => P_HR_S <= "000000101011";
			when "01001101101" => P_HR_S <= "000000100001";
			when "01001101110" => P_HR_S <= "000000100001";
			when "01001101111" => P_HR_S <= "000000001011";
			when "01001110001" => P_HR_S <= "000000100001";
			when "01001110011" => P_HR_S <= "000000010110";
			when "01001110100" => P_HR_S <= "000000010110";
			when "01001110101" => P_HR_S <= "000000001011";
			when "01001110110" => P_HR_S <= "000000101011";
			when "01001111000" => P_HR_S <= "000000010110";
			when "01001111001" => P_HR_S <= "000000100001";
			when "01001111010" => P_HR_S <= "000000100001";
			when "01001111011" => P_HR_S <= "000000010110";
			when "01001111100" => P_HR_S <= "000000001011";
			when "01001111110" => P_HR_S <= "000001100010";
			when "01001111111" => P_HR_S <= "000000101011";
			when "01010000000" => P_HR_S <= "000000101011";
			when "01010000001" => P_HR_S <= "000000110110";
			when "01010000010" => P_HR_S <= "000001000001";
			when "01010000100" => P_HR_S <= "000000100001";
			when "01010000101" => P_HR_S <= "000000101011";
			when "01010000110" => P_HR_S <= "000000101011";
			when "01010001001" => P_HR_S <= "000000110110";
			when "01010001010" => P_HR_S <= "000000100001";
			when "01010001011" => P_HR_S <= "000000010110";
			when "01010001110" => P_HR_S <= "000000010110";
			when "01010001111" => P_HR_S <= "000001000001";
			when "01010010000" => P_HR_S <= "000000001011";
			when "01010010010" => P_HR_S <= "000001010111";
			when "01010010011" => P_HR_S <= "000000010110";
			when "01010010100" => P_HR_S <= "000000010110";
			when "01010010101" => P_HR_S <= "000000010110";
			when "01010010111" => P_HR_S <= "000000001011";
			when "01010011000" => P_HR_S <= "000000100001";
			when "01010011001" => P_HR_S <= "000000100001";
			when "01010011011" => P_HR_S <= "000000110110";
			when "01010011100" => P_HR_S <= "000001000001";
			when "01010011101" => P_HR_S <= "000000010110";
			when "01010011111" => P_HR_S <= "000000101011";
			when "01010100000" => P_HR_S <= "000001000001";
			when "01010100001" => P_HR_S <= "000000100001";
			when "01010100011" => P_HR_S <= "000000100001";
			when "01010100100" => P_HR_S <= "000000010110";
			when "01010100101" => P_HR_S <= "000000001011";
			when "01010100111" => P_HR_S <= "000001001100";
			when "01010101000" => P_HR_S <= "000000010110";
			when "01010101010" => P_HR_S <= "000000010110";
			when "01010101011" => P_HR_S <= "000000010110";
			when "01010101100" => P_HR_S <= "000001000001";
			when "01010101110" => P_HR_S <= "000000110110";
			when "01010101111" => P_HR_S <= "000000100001";
			when "01010110001" => P_HR_S <= "000000010110";
			when "01010110010" => P_HR_S <= "000000100001";
			when "01010110011" => P_HR_S <= "000000010110";
			when "01010110101" => P_HR_S <= "000000100001";
			when "01010110110" => P_HR_S <= "000000101011";
			when "01010111000" => P_HR_S <= "000000010110";
			when "01010111001" => P_HR_S <= "000001000001";
			when "01010111100" => P_HR_S <= "000001001100";
			when "01010111101" => P_HR_S <= "000000100001";
			when "01010111111" => P_HR_S <= "000000110110";
			when "01011000000" => P_HR_S <= "000000010110";
			when "01011000010" => P_HR_S <= "000000010110";
			when "01011000011" => P_HR_S <= "000000100001";
			when "01011000101" => P_HR_S <= "000001001100";
			when "01011000110" => P_HR_S <= "000000100001";
			when "01011001000" => P_HR_S <= "000000101011";
			when "01011001001" => P_HR_S <= "000000010110";
			when "01011001011" => P_HR_S <= "000000010110";
			when "01011001100" => P_HR_S <= "000000100001";
			when "01011001110" => P_HR_S <= "000001010111";
			when "01011001111" => P_HR_S <= "000000110110";
			when "01011010001" => P_HR_S <= "000001000001";
			when "01011010011" => P_HR_S <= "000000010110";
			when "01011010100" => P_HR_S <= "000000101011";
			when "01011010110" => P_HR_S <= "000001001100";
			when "01011010111" => P_HR_S <= "000000101011";
			when "01011011001" => P_HR_S <= "000001000001";
			when "01011011010" => P_HR_S <= "000000101011";
			when "01011011100" => P_HR_S <= "000000010110";
			when "01011011110" => P_HR_S <= "000000110110";
			when "01011011111" => P_HR_S <= "000001000001";
			when "01011100001" => P_HR_S <= "000000110110";
			when "01011100010" => P_HR_S <= "000000100001";
			when "01011100100" => P_HR_S <= "000000100001";
			when "01011100110" => P_HR_S <= "000000101011";
			when "01011100111" => P_HR_S <= "000001010111";
			when "01011101001" => P_HR_S <= "000001000001";
			when "01011101011" => P_HR_S <= "000000101011";
			when "01011101100" => P_HR_S <= "000001000001";
			when "01011101110" => P_HR_S <= "000001001100";
			when "01011110000" => P_HR_S <= "000001000001";
			when "01011110001" => P_HR_S <= "000000001011";
			when "01011110011" => P_HR_S <= "000000100001";
			when "01011110101" => P_HR_S <= "000001000001";
			when "01011110110" => P_HR_S <= "000001000001";
			when "01011111000" => P_HR_S <= "000000100001";
			when "01011111010" => P_HR_S <= "000000110110";
			when "01011111100" => P_HR_S <= "000001000001";
			when "01011111101" => P_HR_S <= "000010000010";
			when "01011111111" => P_HR_S <= "000000010110";
			when "01100000001" => P_HR_S <= "000000101011";
			when "01100000011" => P_HR_S <= "000000001011";
			when "01100000100" => P_HR_S <= "000001001100";
			when "01100000110" => P_HR_S <= "000000101011";
			when "01100001000" => P_HR_S <= "000001100010";
			when "01100001010" => P_HR_S <= "000000010110";
			when "01100001100" => P_HR_S <= "000000101011";
			when "01100001101" => P_HR_S <= "000000110110";
			when "01100001111" => P_HR_S <= "000001010111";
			when "01100010001" => P_HR_S <= "000000100001";
			when "01100010011" => P_HR_S <= "000001010111";
			when "01100010101" => P_HR_S <= "000001000001";
			when "01100010111" => P_HR_S <= "000000100001";
			when "01100011000" => P_HR_S <= "000000110110";
			when "01100011010" => P_HR_S <= "000001001100";
			when "01100011110" => P_HR_S <= "000001001100";
			when "01100100000" => P_HR_S <= "000001100010";
			when "01100100010" => P_HR_S <= "000000010110";
			when "01100100100" => P_HR_S <= "000000001011";
			when "01100100110" => P_HR_S <= "000000100001";
			when "01100101000" => P_HR_S <= "000001101100";
			when "01100101010" => P_HR_S <= "000001100010";
			when "01100101100" => P_HR_S <= "000000100001";
			when "01100101110" => P_HR_S <= "000000001011";
			when "01100110000" => P_HR_S <= "000000010110";
			when "01100110010" => P_HR_S <= "000001000001";
			when "01100110100" => P_HR_S <= "000000100001";
			when "01100110110" => P_HR_S <= "000000101011";
			when "01100111000" => P_HR_S <= "000000100001";
			when "01100111010" => P_HR_S <= "000000110110";
			when "01100111100" => P_HR_S <= "000000100001";
			when "01100111110" => P_HR_S <= "000000110110";
			when "01101000000" => P_HR_S <= "000001000001";
			when "01101000010" => P_HR_S <= "000000101011";
			when "01101000100" => P_HR_S <= "000000101011";
			when "01101000110" => P_HR_S <= "000000001011";
			when "01101001000" => P_HR_S <= "000000010110";
			when "01101001100" => P_HR_S <= "000000100001";
			when "01101001110" => P_HR_S <= "000000110110";
			when "01101010000" => P_HR_S <= "000000001011";
			when "01101010011" => P_HR_S <= "000000110110";
			when "01101010101" => P_HR_S <= "000000010110";
			when "01101010111" => P_HR_S <= "000000001011";
			when "01101011001" => P_HR_S <= "000000001011";
			when "01101011011" => P_HR_S <= "000000101011";
			when "01101011110" => P_HR_S <= "000000001011";
			when "01101100000" => P_HR_S <= "000000100001";
			when "01101100010" => P_HR_S <= "000000001011";
			when "01101100100" => P_HR_S <= "000000101011";
			when "01101100110" => P_HR_S <= "000001000001";
			when "01101101001" => P_HR_S <= "000000100001";
			when "01101101011" => P_HR_S <= "000000001011";
			when "01101101101" => P_HR_S <= "000000010110";
			when "01101110000" => P_HR_S <= "000000001011";
			when "01101110010" => P_HR_S <= "000000010110";
			when "01101110100" => P_HR_S <= "000000010110";
			when "01101111011" => P_HR_S <= "000000010110";
			when "01101111110" => P_HR_S <= "000000001011";
			when "01110000101" => P_HR_S <= "000000001011";
			when "01110000111" => P_HR_S <= "000000010110";
			when "01110001010" => P_HR_S <= "000000010110";
			when "01110001100" => P_HR_S <= "000000010110";
			when "01110001111" => P_HR_S <= "000000010110";
			when "01110010100" => P_HR_S <= "000000010110";
			when "01110010110" => P_HR_S <= "000000001011";
			when "01110011001" => P_HR_S <= "000000001011";
			when "01110011011" => P_HR_S <= "000000001011";
			when "01110100011" => P_HR_S <= "000000001011";
			when "01110101101" => P_HR_S <= "000000001011";
			when "01110110010" => P_HR_S <= "000000010110";
			when "01110110101" => P_HR_S <= "000000001011";
			when "01110111000" => P_HR_S <= "000000100001";
			when "01110111011" => P_HR_S <= "000000001011";
			when "01111000000" => P_HR_S <= "000000001011";
			when "01111000110" => P_HR_S <= "000000001011";
			when "01111001000" => P_HR_S <= "000000001011";
			when "01111001011" => P_HR_S <= "000000010110";
			when "01111001110" => P_HR_S <= "000000010110";
			when "01111010001" => P_HR_S <= "000000010110";
			when "01111010100" => P_HR_S <= "000000010110";
			when "01111010110" => P_HR_S <= "000000001011";
			when "01111011100" => P_HR_S <= "000000001011";
			when "01111011111" => P_HR_S <= "000000001011";
			when "01111100010" => P_HR_S <= "000000001011";
			when "01111100101" => P_HR_S <= "000000010110";
			when "01111101000" => P_HR_S <= "000000001011";
			when "01111101011" => P_HR_S <= "000000100001";
			when "01111101110" => P_HR_S <= "000000010110";
			when "01111110111" => P_HR_S <= "000000100001";
			when "01111111101" => P_HR_S <= "000000101011";
			when "10000000000" => P_HR_S <= "000000001011";
			when "10000000100" => P_HR_S <= "000000001011";
			when "10000000111" => P_HR_S <= "000000010110";
			when "10000001010" => P_HR_S <= "000000100001";
			when "10000001101" => P_HR_S <= "000000001011";
			when "10000010000" => P_HR_S <= "000000101011";
			when "10000010011" => P_HR_S <= "000000100001";
			when "10000010111" => P_HR_S <= "000000100001";
			when "10000011010" => P_HR_S <= "000000101011";
			when "10000011101" => P_HR_S <= "000000101011";
			when "10000100100" => P_HR_S <= "000000010110";
			when "10000101011" => P_HR_S <= "000000100001";
			when "10000101110" => P_HR_S <= "000000010110";
			when "10000110001" => P_HR_S <= "000000001011";
			when "10000111000" => P_HR_S <= "000000001011";
			when others        => P_HR_S <= "000000000001";
		end case;
		
        --stress_score_temp <= P_TEMP_S * P_STRESS * P_EDA_S * P_HR_S;
        --stress_score_temp <= P_TEMP_S * P_EDA_S * P_HR_S;
	end process;
	
	process(P_TEMP_S,P_EDA_S,P_HR_S)
	begin
	stress_score_temp <= P_TEMP_S * P_STRESS * P_EDA_S * P_HR_S;
	end process;
	
	process(P_TEMP_NS,P_EDA_NS,P_HR_NS)
	begin
	not_stress_score_temp <= P_TEMP_NS * P_NOT_STRESS * P_EDA_NS * P_HR_NS;
	end process;
	
	process(temp, eda, hr)
	begin
		case temp is
			when "011110110" => P_TEMP_NS <= "000010110000";
			when "011110111" => P_TEMP_NS <= "001100101110";
			when "011111000" => P_TEMP_NS <= "001000001111";
			when "011111001" => P_TEMP_NS <= "000001111100";
			when "011111010" => P_TEMP_NS <= "000110011100";
			when "011111011" => P_TEMP_NS <= "000111010000";
			when "011111100" => P_TEMP_NS <= "001000100011";
			when "011111101" => P_TEMP_NS <= "001100101010";
			when "011111110" => P_TEMP_NS <= "000011110000";
			when "011111111" => P_TEMP_NS <= "000011000011";
			when "100000000" => P_TEMP_NS <= "000100001010";
			when "100000001" => P_TEMP_NS <= "000000101111";
			when "100000010" => P_TEMP_NS <= "000000110110";
			when "100000011" => P_TEMP_NS <= "000000100101";
			when "100000100" => P_TEMP_NS <= "000011010001";
			when "100000101" => P_TEMP_NS <= "000001101011";
			when "100000110" => P_TEMP_NS <= "000000101110";
			when "100000111" => P_TEMP_NS <= "001001001001";
			when "100001000" => P_TEMP_NS <= "010000100100";
			when "100001001" => P_TEMP_NS <= "010101101000";
			when "100001010" => P_TEMP_NS <= "001101100101";
			when "100001011" => P_TEMP_NS <= "001111111010";
			when "100001100" => P_TEMP_NS <= "000000000111";
			when others      => P_TEMP_NS <= "000000000001";
		end case;	
	
		case hr is
			when "00100010111" => P_HR_NS <= "000000000100";
			when "00100011111" => P_HR_NS <= "000000000100";
			when "00100100001" => P_HR_NS <= "000000000100";
			when "00100101010" => P_HR_NS <= "000000001001";
			when "00100101011" => P_HR_NS <= "000000000100";
			when "00100110000" => P_HR_NS <= "000000000100";
			when "00100110011" => P_HR_NS <= "000000001001";
			when "00100110110" => P_HR_NS <= "000000001001";
			when "00100111000" => P_HR_NS <= "000000000100";
			when "00100111010" => P_HR_NS <= "000000000100";
			when "00100111011" => P_HR_NS <= "000000001001";
			when "00100111110" => P_HR_NS <= "000000001001";
			when "00100111111" => P_HR_NS <= "000000000100";
			when "00101000000" => P_HR_NS <= "000000001101";
			when "00101000010" => P_HR_NS <= "000000001001";
			when "00101000011" => P_HR_NS <= "000000001001";
			when "00101000100" => P_HR_NS <= "000000000100";
			when "00101000101" => P_HR_NS <= "000000000100";
			when "00101000110" => P_HR_NS <= "000000001001";
			when "00101000111" => P_HR_NS <= "000000001001";
			when "00101001000" => P_HR_NS <= "000000001001";
			when "00101001011" => P_HR_NS <= "000000001101";
			when "00101001110" => P_HR_NS <= "000000000100";
			when "00101001111" => P_HR_NS <= "000000001001";
			when "00101010000" => P_HR_NS <= "000000000100";
			when "00101010001" => P_HR_NS <= "000000010010";
			when "00101010010" => P_HR_NS <= "000000010010";
			when "00101010100" => P_HR_NS <= "000000011011";
			when "00101010101" => P_HR_NS <= "000000001001";
			when "00101010110" => P_HR_NS <= "000000001001";
			when "00101010111" => P_HR_NS <= "000000010010";
			when "00101011000" => P_HR_NS <= "000000010110";
			when "00101011001" => P_HR_NS <= "000000001001";
			when "00101011010" => P_HR_NS <= "000000010110";
			when "00101011011" => P_HR_NS <= "000000010010";
			when "00101011100" => P_HR_NS <= "000000001001";
			when "00101011101" => P_HR_NS <= "000000011011";
			when "00101011110" => P_HR_NS <= "000000001101";
			when "00101011111" => P_HR_NS <= "000000000100";
			when "00101100000" => P_HR_NS <= "000000001001";
			when "00101100001" => P_HR_NS <= "000000010010";
			when "00101100010" => P_HR_NS <= "000000010110";
			when "00101100011" => P_HR_NS <= "000000010010";
			when "00101100100" => P_HR_NS <= "000000010110";
			when "00101100101" => P_HR_NS <= "000000011111";
			when "00101100110" => P_HR_NS <= "000000000100";
			when "00101100111" => P_HR_NS <= "000000101101";
			when "00101101000" => P_HR_NS <= "000000011011";
			when "00101101001" => P_HR_NS <= "000000101101";
			when "00101101010" => P_HR_NS <= "000000110001";
			when "00101101011" => P_HR_NS <= "000000011111";
			when "00101101100" => P_HR_NS <= "000000011111";
			when "00101101101" => P_HR_NS <= "000000100100";
			when "00101101110" => P_HR_NS <= "000001001100";
			when "00101101111" => P_HR_NS <= "000000101101";
			when "00101110000" => P_HR_NS <= "000000111110";
			when "00101110001" => P_HR_NS <= "000000011111";
			when "00101110010" => P_HR_NS <= "000001001100";
			when "00101110011" => P_HR_NS <= "000000101000";
			when "00101110100" => P_HR_NS <= "000000011011";
			when "00101110101" => P_HR_NS <= "000000100100";
			when "00101110110" => P_HR_NS <= "000000100100";
			when "00101110111" => P_HR_NS <= "000001001100";
			when "00101111000" => P_HR_NS <= "000001000111";
			when "00101111001" => P_HR_NS <= "000000101101";
			when "00101111010" => P_HR_NS <= "000000110001";
			when "00101111011" => P_HR_NS <= "000000101000";
			when "00101111100" => P_HR_NS <= "000000011011";
			when "00101111101" => P_HR_NS <= "000001011001";
			when "00101111110" => P_HR_NS <= "000000110001";
			when "00101111111" => P_HR_NS <= "000000010110";
			when "00110000000" => P_HR_NS <= "000001010101";
			when "00110000001" => P_HR_NS <= "000000100100";
			when "00110000010" => P_HR_NS <= "000000011011";
			when "00110000011" => P_HR_NS <= "000001000011";
			when "00110000100" => P_HR_NS <= "000001101111";
			when "00110000101" => P_HR_NS <= "000000101101";
			when "00110000110" => P_HR_NS <= "000001000011";
			when "00110000111" => P_HR_NS <= "000001001100";
			when "00110001000" => P_HR_NS <= "000000110001";
			when "00110001001" => P_HR_NS <= "000010001010";
			when "00110001010" => P_HR_NS <= "000000111110";
			when "00110001011" => P_HR_NS <= "000001000011";
			when "00110001100" => P_HR_NS <= "000001011001";
			when "00110001101" => P_HR_NS <= "000000111110";
			when "00110001110" => P_HR_NS <= "000001011101";
			when "00110001111" => P_HR_NS <= "000000101101";
			when "00110010000" => P_HR_NS <= "000010001110";
			when "00110010001" => P_HR_NS <= "000001011001";
			when "00110010010" => P_HR_NS <= "000001100110";
			when "00110010011" => P_HR_NS <= "000001100010";
			when "00110010100" => P_HR_NS <= "000001001100";
			when "00110010101" => P_HR_NS <= "000001010101";
			when "00110010110" => P_HR_NS <= "000001010101";
			when "00110010111" => P_HR_NS <= "000001111101";
			when "00110011000" => P_HR_NS <= "000001100010";
			when "00110011001" => P_HR_NS <= "000001100010";
			when "00110011010" => P_HR_NS <= "000001110100";
			when "00110011011" => P_HR_NS <= "000000111110";
			when "00110011100" => P_HR_NS <= "000001010000";
			when "00110011101" => P_HR_NS <= "000000111110";
			when "00110011110" => P_HR_NS <= "000001010000";
			when "00110011111" => P_HR_NS <= "000000110101";
			when "00110100000" => P_HR_NS <= "000001011001";
			when "00110100001" => P_HR_NS <= "000001010101";
			when "00110100010" => P_HR_NS <= "000001010000";
			when "00110100011" => P_HR_NS <= "000000110101";
			when "00110100100" => P_HR_NS <= "000000101101";
			when "00110100101" => P_HR_NS <= "000001000011";
			when "00110100110" => P_HR_NS <= "000001010101";
			when "00110100111" => P_HR_NS <= "000001000011";
			when "00110101000" => P_HR_NS <= "000000111010";
			when "00110101001" => P_HR_NS <= "000001000011";
			when "00110101010" => P_HR_NS <= "000001100110";
			when "00110101011" => P_HR_NS <= "000000111010";
			when "00110101100" => P_HR_NS <= "000000110101";
			when "00110101101" => P_HR_NS <= "000001011001";
			when "00110101110" => P_HR_NS <= "000000110001";
			when "00110101111" => P_HR_NS <= "000000101101";
			when "00110110000" => P_HR_NS <= "000001011001";
			when "00110110001" => P_HR_NS <= "000000011011";
			when "00110110010" => P_HR_NS <= "000001010101";
			when "00110110011" => P_HR_NS <= "000001000111";
			when "00110110100" => P_HR_NS <= "000001100010";
			when "00110110101" => P_HR_NS <= "000000110101";
			when "00110110110" => P_HR_NS <= "000000111010";
			when "00110110111" => P_HR_NS <= "000000110101";
			when "00110111000" => P_HR_NS <= "000001000011";
			when "00110111001" => P_HR_NS <= "000000011011";
			when "00110111010" => P_HR_NS <= "000000111110";
			when "00110111011" => P_HR_NS <= "000001010000";
			when "00110111100" => P_HR_NS <= "000000111010";
			when "00110111101" => P_HR_NS <= "000000101000";
			when "00110111110" => P_HR_NS <= "000000101000";
			when "00110111111" => P_HR_NS <= "000000111110";
			when "00111000000" => P_HR_NS <= "000000110001";
			when "00111000001" => P_HR_NS <= "000001000011";
			when "00111000010" => P_HR_NS <= "000001000111";
			when "00111000011" => P_HR_NS <= "000000010010";
			when "00111000100" => P_HR_NS <= "000000101101";
			when "00111000101" => P_HR_NS <= "000000110101";
			when "00111000110" => P_HR_NS <= "000000100100";
			when "00111000111" => P_HR_NS <= "000000010110";
			when "00111001000" => P_HR_NS <= "000000010110";
			when "00111001001" => P_HR_NS <= "000000111010";
			when "00111001010" => P_HR_NS <= "000000111010";
			when "00111001011" => P_HR_NS <= "000000010010";
			when "00111001100" => P_HR_NS <= "000000110001";
			when "00111001101" => P_HR_NS <= "000000011011";
			when "00111001110" => P_HR_NS <= "000000110001";
			when "00111001111" => P_HR_NS <= "000000101000";
			when "00111010000" => P_HR_NS <= "000000001001";
			when "00111010001" => P_HR_NS <= "000000011111";
			when "00111010010" => P_HR_NS <= "000000011011";
			when "00111010011" => P_HR_NS <= "000001001100";
			when "00111010100" => P_HR_NS <= "000000100100";
			when "00111010101" => P_HR_NS <= "000000111110";
			when "00111010110" => P_HR_NS <= "000000100100";
			when "00111010111" => P_HR_NS <= "000000111010";
			when "00111011000" => P_HR_NS <= "000000101000";
			when "00111011001" => P_HR_NS <= "000001000111";
			when "00111011010" => P_HR_NS <= "000000011111";
			when "00111011011" => P_HR_NS <= "000000011011";
			when "00111011100" => P_HR_NS <= "000000101000";
			when "00111011101" => P_HR_NS <= "000000101101";
			when "00111011110" => P_HR_NS <= "000000100100";
			when "00111011111" => P_HR_NS <= "000001001100";
			when "00111100000" => P_HR_NS <= "000000011111";
			when "00111100001" => P_HR_NS <= "000000100100";
			when "00111100010" => P_HR_NS <= "000000001001";
			when "00111100011" => P_HR_NS <= "000000011011";
			when "00111100100" => P_HR_NS <= "000000001001";
			when "00111100101" => P_HR_NS <= "000000101101";
			when "00111100110" => P_HR_NS <= "000001000011";
			when "00111100111" => P_HR_NS <= "000000010110";
			when "00111101000" => P_HR_NS <= "000000011111";
			when "00111101001" => P_HR_NS <= "000000010010";
			when "00111101010" => P_HR_NS <= "000000010010";
			when "00111101011" => P_HR_NS <= "000000010110";
			when "00111101100" => P_HR_NS <= "000000010110";
			when "00111101101" => P_HR_NS <= "000000010110";
			when "00111101111" => P_HR_NS <= "000000101000";
			when "00111110000" => P_HR_NS <= "000000101000";
			when "00111110001" => P_HR_NS <= "000000001001";
			when "00111110010" => P_HR_NS <= "000000010010";
			when "00111110011" => P_HR_NS <= "000000101101";
			when "00111110100" => P_HR_NS <= "000000010010";
			when "00111110101" => P_HR_NS <= "000000010110";
			when "00111110110" => P_HR_NS <= "000000000100";
			when "00111110111" => P_HR_NS <= "000000010010";
			when "00111111000" => P_HR_NS <= "000000001101";
			when "00111111001" => P_HR_NS <= "000000101101";
			when "00111111010" => P_HR_NS <= "000000001101";
			when "00111111011" => P_HR_NS <= "000000011011";
			when "00111111100" => P_HR_NS <= "000000011111";
			when "00111111101" => P_HR_NS <= "000000010010";
			when "00111111110" => P_HR_NS <= "000000011011";
			when "00111111111" => P_HR_NS <= "000000010110";
			when "01000000000" => P_HR_NS <= "000000010010";
			when "01000000001" => P_HR_NS <= "000000001001";
			when "01000000010" => P_HR_NS <= "000000010010";
			when "01000000011" => P_HR_NS <= "000000101101";
			when "01000000100" => P_HR_NS <= "000000011011";
			when "01000000101" => P_HR_NS <= "000000001101";
			when "01000000110" => P_HR_NS <= "000000010010";
			when "01000000111" => P_HR_NS <= "000000110101";
			when "01000001000" => P_HR_NS <= "000000001101";
			when "01000001001" => P_HR_NS <= "000000001101";
			when "01000001010" => P_HR_NS <= "000000001101";
			when "01000001011" => P_HR_NS <= "000000100100";
			when "01000001100" => P_HR_NS <= "000000011011";
			when "01000001101" => P_HR_NS <= "000000000100";
			when "01000001110" => P_HR_NS <= "000000010010";
			when "01000001111" => P_HR_NS <= "000000100100";
			when "01000010000" => P_HR_NS <= "000000001101";
			when "01000010001" => P_HR_NS <= "000000001001";
			when "01000010010" => P_HR_NS <= "000000011011";
			when "01000010011" => P_HR_NS <= "000000011011";
			when "01000010100" => P_HR_NS <= "000000110001";
			when "01000010101" => P_HR_NS <= "000000010010";
			when "01000010110" => P_HR_NS <= "000000011111";
			when "01000010111" => P_HR_NS <= "000000001101";
			when "01000011000" => P_HR_NS <= "000000011111";
			when "01000011001" => P_HR_NS <= "000000010010";
			when "01000011010" => P_HR_NS <= "000000001001";
			when "01000011011" => P_HR_NS <= "000000001101";
			when "01000011100" => P_HR_NS <= "000000011111";
			when "01000011101" => P_HR_NS <= "000000001001";
			when "01000011110" => P_HR_NS <= "000000001101";
			when "01000011111" => P_HR_NS <= "000000001101";
			when "01000100000" => P_HR_NS <= "000000100100";
			when "01000100001" => P_HR_NS <= "000000010110";
			when "01000100010" => P_HR_NS <= "000000001101";
			when "01000100011" => P_HR_NS <= "000000001101";
			when "01000100100" => P_HR_NS <= "000000010110";
			when "01000100101" => P_HR_NS <= "000000010010";
			when "01000100110" => P_HR_NS <= "000000010110";
			when "01000100111" => P_HR_NS <= "000000010010";
			when "01000101000" => P_HR_NS <= "000000001001";
			when "01000101001" => P_HR_NS <= "000000000100";
			when "01000101010" => P_HR_NS <= "000000011011";
			when "01000101011" => P_HR_NS <= "000000010010";
			when "01000101100" => P_HR_NS <= "000000001001";
			when "01000101101" => P_HR_NS <= "000000001001";
			when "01000101110" => P_HR_NS <= "000000011011";
			when "01000101111" => P_HR_NS <= "000000001101";
			when "01000110000" => P_HR_NS <= "000000001001";
			when "01000110001" => P_HR_NS <= "000000010110";
			when "01000110010" => P_HR_NS <= "000000001101";
			when "01000110011" => P_HR_NS <= "000000000100";
			when "01000110100" => P_HR_NS <= "000000001001";
			when "01000110110" => P_HR_NS <= "000000001101";
			when "01000110111" => P_HR_NS <= "000000001001";
			when "01000111000" => P_HR_NS <= "000000001101";
			when "01000111001" => P_HR_NS <= "000000011011";
			when "01000111010" => P_HR_NS <= "000000000100";
			when "01000111011" => P_HR_NS <= "000000001101";
			when "01000111100" => P_HR_NS <= "000000010110";
			when "01000111101" => P_HR_NS <= "000000001001";
			when "01000111110" => P_HR_NS <= "000000001001";
			when "01000111111" => P_HR_NS <= "000000010010";
			when "01001000001" => P_HR_NS <= "000000001001";
			when "01001000010" => P_HR_NS <= "000000001101";
			when "01001000011" => P_HR_NS <= "000000001101";
			when "01001000100" => P_HR_NS <= "000000000100";
			when "01001000101" => P_HR_NS <= "000000000100";
			when "01001000110" => P_HR_NS <= "000000010110";
			when "01001000111" => P_HR_NS <= "000000001101";
			when "01001001000" => P_HR_NS <= "000000010110";
			when "01001001001" => P_HR_NS <= "000000010010";
			when "01001001010" => P_HR_NS <= "000000000100";
			when "01001001011" => P_HR_NS <= "000000001001";
			when "01001001100" => P_HR_NS <= "000000000100";
			when "01001001101" => P_HR_NS <= "000000001101";
			when "01001001111" => P_HR_NS <= "000000000100";
			when "01001010000" => P_HR_NS <= "000000000100";
			when "01001010001" => P_HR_NS <= "000000001001";
			when "01001010010" => P_HR_NS <= "000000000100";
			when "01001010100" => P_HR_NS <= "000000000100";
			when "01001010101" => P_HR_NS <= "000000001001";
			when "01001010110" => P_HR_NS <= "000000001001";
			when "01001010111" => P_HR_NS <= "000000000100";
			when "01001011000" => P_HR_NS <= "000000001101";
			when "01001011001" => P_HR_NS <= "000000001101";
			when "01001011010" => P_HR_NS <= "000000000100";
			when "01001011011" => P_HR_NS <= "000000000100";
			when "01001011101" => P_HR_NS <= "000000000100";
			when "01001011110" => P_HR_NS <= "000000000100";
			when "01001100000" => P_HR_NS <= "000000000100";
			when "01001100010" => P_HR_NS <= "000000001001";
			when "01001100011" => P_HR_NS <= "000000000100";
			when "01001100101" => P_HR_NS <= "000000001001";
			when "01001100110" => P_HR_NS <= "000000001101";
			when "01001100111" => P_HR_NS <= "000000000100";
			when "01001101001" => P_HR_NS <= "000000000100";
			when "01001101010" => P_HR_NS <= "000000000100";
			when "01001101100" => P_HR_NS <= "000000000100";
			when "01001101110" => P_HR_NS <= "000000000100";
			when "01001101111" => P_HR_NS <= "000000000100";
			when "01010000000" => P_HR_NS <= "000000000100";
			when "01010000001" => P_HR_NS <= "000000000100";
			when "01010000100" => P_HR_NS <= "000000000100";
			when "01010000110" => P_HR_NS <= "000000000100";
			when "01010001001" => P_HR_NS <= "000000000100";
			when "01010001010" => P_HR_NS <= "000000000100";
			when "01010011111" => P_HR_NS <= "000000000100";
			when "01010100101" => P_HR_NS <= "000000000100";
			when "01010101000" => P_HR_NS <= "000000000100";
			when "01010101010" => P_HR_NS <= "000000000100";
			when others       => P_HR_NS <= "000000000001";
		end case;

		case eda is
			when "0110100" => P_EDA_NS <= "000000111110";
			when "0110101" => P_EDA_NS <= "000111000011";
			when "0110110" => P_EDA_NS <= "001001001000";
			when "0110111" => P_EDA_NS <= "000010110010";
			when "0111000" => P_EDA_NS <= "000101001000";
			when "0111001" => P_EDA_NS <= "001110010000";
			when "0111010" => P_EDA_NS <= "001010010111";
			when "0111011" => P_EDA_NS <= "001001001001";
			when "0111100" => P_EDA_NS <= "001001111001";
			when "0111101" => P_EDA_NS <= "000001111000";
			when "0111110" => P_EDA_NS <= "000110000110";
			when "0111111" => P_EDA_NS <= "000111111000";
			when "0100000" => P_EDA_NS <= "000101101101";
			when "1000001" => P_EDA_NS <= "000110111001";
            when "1000010" => P_EDA_NS <= "000101100011";
            when "1000011" => P_EDA_NS <= "000000101100";
            when "1000100" => P_EDA_NS <= "000000111110";
            when "1000101" => P_EDA_NS <= "000001001000";
            when "1000110" => P_EDA_NS <= "000010010101";
            when "1000111" => P_EDA_NS <= "000000011110";
			when others   => P_EDA_NS <= "000000000001";
		end case;
		
		--not_stress_score_temp <= P_TEMP_NS * P_NOT_STRESS * P_EDA_NS * P_HR_NS;
		--not_stress_score_temp <= ('0'&P_TEMP_NS) * P_NOT_STRESS * ('0'&P_EDA_NS) * ('0'&P_HR_NS);
	end process;
	
	process(clk, rst)
	begin
		if (rst = '1') then
			stress_score <= (others => '0');
			not_stress_score <= (others => '0');
			status <= (others => '0');
		elsif (rising_edge(clk)) then
		
			stress_score <= std_logic_vector(stress_score_temp);
			not_stress_score <= std_logic_vector(not_stress_score_temp);
			
		    if stress_score_temp < not_stress_score_temp then
		        status <= "01"; -- not stressed
			elsif stress_score_temp > not_stress_score_temp then
				status <= "10"; -- stressed
			elsif stress_score_temp = not_stress_score_temp then
				status <= "11"; -- rare, equality
			else
				status <= "00";
			end if;
		end if;
	end process;

end behavioral;