-----------------------------------------------------------------
-- Created By: Richard Cho
-- Create Date: 3/17/2022
-----------------------------------------------------------------
-- Naive Bayes model for stress detection using the WESAD
-- database. Training mode increases individual probability
-- values based on given inputs.
-- Two machines run in parallel to calculate a stress and
-- non-stress score. Whichever score is higher is the final
-- decision. If scores are equal (highly unlikely) then it
-- should choose not stressed as the default (not in yet).
-----------------------------------------------------------------
-- Revision History
-- 3/17/2022: Created model for S2 only
-- 4/24/2022: Updated model for S2 and S3 combined
-- 5/28/22: Updated model for every WESAD subject
-----------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity SCORE_CALC_T is
    
    port (
        clk : in std_logic; -- system clock
        rst : in std_logic; -- system reset
		temp : in std_logic_vector (8 downto 0); -- celcius
		eda : in std_logic_vector (7 downto 0); --micro siemens
		hr : in std_logic_vector (10 downto 0); -- bpm
		s1 : in std_logic_vector (1 downto 0); -- switch for states
		status : out std_logic_vector (1 downto 0)); -- output
		
end SCORE_CALC_T;

architecture behavioral of SCORE_CALC_T is
	
	signal P_TEMP_S1 : unsigned(11 downto 0);
	signal P_TEMP_S2 : unsigned(11 downto 0);
	signal P_TEMP_S3 : unsigned(11 downto 0);
	signal P_TEMP_S4 : unsigned(11 downto 0);
	signal P_TEMP_S5 : unsigned(11 downto 0);
	signal P_TEMP_S6 : unsigned(11 downto 0);
	signal P_TEMP_S7 : unsigned(11 downto 0);
	signal P_TEMP_S8 : unsigned(11 downto 0);
	signal P_TEMP_S9 : unsigned(11 downto 0);
	signal P_TEMP_S10 : unsigned(11 downto 0);
	signal P_TEMP_S11 : unsigned(11 downto 0);
	signal P_TEMP_S12 : unsigned(11 downto 0);
	signal P_TEMP_S13 : unsigned(11 downto 0);
	signal P_TEMP_S14 : unsigned(11 downto 0);
	signal P_TEMP_S15 : unsigned(11 downto 0);
	signal P_TEMP_S16 : unsigned(11 downto 0);
	signal P_TEMP_S17 : unsigned(11 downto 0);
	signal P_TEMP_S18 : unsigned(11 downto 0);
	signal P_TEMP_S19 : unsigned(11 downto 0);
	signal P_TEMP_S20 : unsigned(11 downto 0);
	signal P_TEMP_S21 : unsigned(11 downto 0);
	signal P_TEMP_S22 : unsigned(11 downto 0);
	signal P_TEMP_S23 : unsigned(11 downto 0);
	signal P_TEMP_S24 : unsigned(11 downto 0);
	signal P_TEMP_S25 : unsigned(11 downto 0);
	signal P_TEMP_S26 : unsigned(11 downto 0);
	signal P_TEMP_S27 : unsigned(11 downto 0);
	signal P_TEMP_S28 : unsigned(11 downto 0);
	signal P_TEMP_S29 : unsigned(11 downto 0);
	signal P_TEMP_S30 : unsigned(11 downto 0);
	signal P_TEMP_S31 : unsigned(11 downto 0);
	signal P_TEMP_S32 : unsigned(11 downto 0);
	signal P_TEMP_S33 : unsigned(11 downto 0);
	signal P_TEMP_S34 : unsigned(11 downto 0);
	signal P_TEMP_S35 : unsigned(11 downto 0);
	signal P_TEMP_S36 : unsigned(11 downto 0);
	signal P_TEMP_S37 : unsigned(11 downto 0);
	signal P_TEMP_S38 : unsigned(11 downto 0);
	signal P_TEMP_S39 : unsigned(11 downto 0);
	signal P_TEMP_S40 : unsigned(11 downto 0);
	

	signal P_EDA_S1 : unsigned(11 downto 0);
	signal P_EDA_S2 : unsigned(11 downto 0);
	signal P_EDA_S3 : unsigned(11 downto 0);
	signal P_EDA_S4 : unsigned(11 downto 0);
	signal P_EDA_S5 : unsigned(11 downto 0);
	signal P_EDA_S6 : unsigned(11 downto 0);
	signal P_EDA_S7 : unsigned(11 downto 0);
	signal P_EDA_S8 : unsigned(11 downto 0);
	signal P_EDA_S9 : unsigned(11 downto 0);
	signal P_EDA_S10 : unsigned(11 downto 0);
	signal P_EDA_S11 : unsigned(11 downto 0);
	signal P_EDA_S12 : unsigned(11 downto 0);
	signal P_EDA_S13 : unsigned(11 downto 0);
	signal P_EDA_S14 : unsigned(11 downto 0);
	signal P_EDA_S15 : unsigned(11 downto 0);
	signal P_EDA_S16 : unsigned(11 downto 0);
	signal P_EDA_S17 : unsigned(11 downto 0);
	signal P_EDA_S18 : unsigned(11 downto 0);
	signal P_EDA_S19 : unsigned(11 downto 0);
	signal P_EDA_S20 : unsigned(11 downto 0);
	signal P_EDA_S21 : unsigned(11 downto 0);
	signal P_EDA_S22 : unsigned(11 downto 0);
	signal P_EDA_S23 : unsigned(11 downto 0);
	signal P_EDA_S24 : unsigned(11 downto 0);
	signal P_EDA_S25 : unsigned(11 downto 0);
	signal P_EDA_S26 : unsigned(11 downto 0);
	signal P_EDA_S27 : unsigned(11 downto 0);
	signal P_EDA_S28 : unsigned(11 downto 0);
	signal P_EDA_S29 : unsigned(11 downto 0);
	signal P_EDA_S30 : unsigned(11 downto 0);
	signal P_EDA_S31 : unsigned(11 downto 0);
	signal P_EDA_S32 : unsigned(11 downto 0);
	signal P_EDA_S33 : unsigned(11 downto 0);
	signal P_EDA_S34 : unsigned(11 downto 0);
	signal P_EDA_S35 : unsigned(11 downto 0);
	signal P_EDA_S36 : unsigned(11 downto 0);
	signal P_EDA_S37 : unsigned(11 downto 0);
	signal P_EDA_S38 : unsigned(11 downto 0);
	signal P_EDA_S39 : unsigned(11 downto 0);
	signal P_EDA_S40 : unsigned(11 downto 0);
	signal P_EDA_S41 : unsigned(11 downto 0);
	signal P_EDA_S42 : unsigned(11 downto 0);
	signal P_EDA_S43 : unsigned(11 downto 0);
	signal P_EDA_S44 : unsigned(11 downto 0);
	signal P_EDA_S45 : unsigned(11 downto 0);
	signal P_EDA_S46 : unsigned(11 downto 0);
	signal P_EDA_S47 : unsigned(11 downto 0);
	signal P_EDA_S48 : unsigned(11 downto 0);
	signal P_EDA_S49 : unsigned(11 downto 0);
	signal P_EDA_S50 : unsigned(11 downto 0);
	signal P_EDA_S51 : unsigned(11 downto 0);
	signal P_EDA_S52 : unsigned(11 downto 0);
	signal P_EDA_S53 : unsigned(11 downto 0);
	signal P_EDA_S54 : unsigned(11 downto 0);
	signal P_EDA_S55 : unsigned(11 downto 0);
	signal P_EDA_S56 : unsigned(11 downto 0);
	signal P_EDA_S57 : unsigned(11 downto 0);
	signal P_EDA_S58 : unsigned(11 downto 0);
	signal P_EDA_S59 : unsigned(11 downto 0);
	signal P_EDA_S60 : unsigned(11 downto 0);
	signal P_EDA_S61 : unsigned(11 downto 0);
	signal P_EDA_S62 : unsigned(11 downto 0);
	signal P_EDA_S63 : unsigned(11 downto 0);
	signal P_EDA_S64 : unsigned(11 downto 0);
	signal P_EDA_S65 : unsigned(11 downto 0);
	signal P_EDA_S66 : unsigned(11 downto 0);
	signal P_EDA_S67 : unsigned(11 downto 0);
	signal P_EDA_S68 : unsigned(11 downto 0);
	signal P_EDA_S69 : unsigned(11 downto 0);
	signal P_EDA_S70 : unsigned(11 downto 0);
	signal P_EDA_S71 : unsigned(11 downto 0);
	signal P_EDA_S72 : unsigned(11 downto 0);
	signal P_EDA_S73 : unsigned(11 downto 0);
	signal P_EDA_S74 : unsigned(11 downto 0);
	signal P_EDA_S75 : unsigned(11 downto 0);
	signal P_EDA_S76 : unsigned(11 downto 0);
	signal P_EDA_S77 : unsigned(11 downto 0);
	signal P_EDA_S78 : unsigned(11 downto 0);
	signal P_EDA_S79 : unsigned(11 downto 0);
	signal P_EDA_S80 : unsigned(11 downto 0);
	signal P_EDA_S81 : unsigned(11 downto 0);
	signal P_EDA_S82 : unsigned(11 downto 0);
	signal P_EDA_S83 : unsigned(11 downto 0);
	signal P_EDA_S84 : unsigned(11 downto 0);
	signal P_EDA_S85 : unsigned(11 downto 0);
	signal P_EDA_S86 : unsigned(11 downto 0);
	signal P_EDA_S87 : unsigned(11 downto 0);
	signal P_EDA_S88 : unsigned(11 downto 0);
	signal P_EDA_S89 : unsigned(11 downto 0);
	signal P_EDA_S90 : unsigned(11 downto 0);
	signal P_EDA_S91 : unsigned(11 downto 0);
	signal P_EDA_S92 : unsigned(11 downto 0);
	signal P_EDA_S93 : unsigned(11 downto 0);
	signal P_EDA_S94 : unsigned(11 downto 0);
	signal P_EDA_S95 : unsigned(11 downto 0);
	signal P_EDA_S96 : unsigned(11 downto 0);
	signal P_EDA_S97 : unsigned(11 downto 0);
	signal P_EDA_S98 : unsigned(11 downto 0);
	signal P_EDA_S99 : unsigned(11 downto 0);
	signal P_EDA_S100 : unsigned(11 downto 0);
	signal P_EDA_S101 : unsigned(11 downto 0);
	signal P_EDA_S102 : unsigned(11 downto 0);
	signal P_EDA_S103 : unsigned(11 downto 0);
	signal P_EDA_S104 : unsigned(11 downto 0);
	signal P_EDA_S105 : unsigned(11 downto 0);
	signal P_EDA_S106 : unsigned(11 downto 0);
	signal P_EDA_S107 : unsigned(11 downto 0);
	signal P_EDA_S108 : unsigned(11 downto 0);
	signal P_EDA_S109 : unsigned(11 downto 0);
	signal P_EDA_S110 : unsigned(11 downto 0);
	signal P_EDA_S111 : unsigned(11 downto 0);
	signal P_EDA_S112 : unsigned(11 downto 0);
	signal P_EDA_S113 : unsigned(11 downto 0);
	signal P_EDA_S114 : unsigned(11 downto 0);
	signal P_EDA_S115 : unsigned(11 downto 0);
	signal P_EDA_S116 : unsigned(11 downto 0);
	signal P_EDA_S117 : unsigned(11 downto 0);
	signal P_EDA_S118 : unsigned(11 downto 0);
	signal P_EDA_S119 : unsigned(11 downto 0);
	signal P_EDA_S120 : unsigned(11 downto 0);
	signal P_EDA_S121 : unsigned(11 downto 0);
	signal P_EDA_S122 : unsigned(11 downto 0);
	signal P_EDA_S123 : unsigned(11 downto 0);
	signal P_EDA_S124 : unsigned(11 downto 0);
	signal P_EDA_S125 : unsigned(11 downto 0);
	signal P_EDA_S126 : unsigned(11 downto 0);
	signal P_EDA_S127 : unsigned(11 downto 0);
	signal P_EDA_S128 : unsigned(11 downto 0);
	signal P_EDA_S129 : unsigned(11 downto 0);
	signal P_EDA_S130 : unsigned(11 downto 0);
	
	signal P_HR_S1 : unsigned(11 downto 0); 
	signal P_HR_S2 : unsigned(11 downto 0); 
	signal P_HR_S3 : unsigned(11 downto 0); 
	signal P_HR_S4 : unsigned(11 downto 0); 
	signal P_HR_S5 : unsigned(11 downto 0); 
	signal P_HR_S6 : unsigned(11 downto 0); 
	signal P_HR_S7 : unsigned(11 downto 0); 
	signal P_HR_S8 : unsigned(11 downto 0); 
	signal P_HR_S9 : unsigned(11 downto 0); 
	signal P_HR_S10 : unsigned(11 downto 0);
	signal P_HR_S11 : unsigned(11 downto 0);
	signal P_HR_S12 : unsigned(11 downto 0);
	signal P_HR_S13 : unsigned(11 downto 0);
	signal P_HR_S14 : unsigned(11 downto 0);
	signal P_HR_S15 : unsigned(11 downto 0);
	signal P_HR_S16 : unsigned(11 downto 0);
	signal P_HR_S17 : unsigned(11 downto 0);
	signal P_HR_S18 : unsigned(11 downto 0);
	signal P_HR_S19 : unsigned(11 downto 0);
	signal P_HR_S20 : unsigned(11 downto 0);
	signal P_HR_S21 : unsigned(11 downto 0);
	signal P_HR_S22 : unsigned(11 downto 0);
	signal P_HR_S23 : unsigned(11 downto 0);
	signal P_HR_S24 : unsigned(11 downto 0);
	signal P_HR_S25 : unsigned(11 downto 0);
	signal P_HR_S26 : unsigned(11 downto 0);
	signal P_HR_S27 : unsigned(11 downto 0);
	signal P_HR_S28 : unsigned(11 downto 0);
	signal P_HR_S29 : unsigned(11 downto 0);
	signal P_HR_S30 : unsigned(11 downto 0);
	signal P_HR_S31 : unsigned(11 downto 0);
	signal P_HR_S32 : unsigned(11 downto 0);
	signal P_HR_S33 : unsigned(11 downto 0);
	signal P_HR_S34 : unsigned(11 downto 0);
	signal P_HR_S35 : unsigned(11 downto 0);
	signal P_HR_S36 : unsigned(11 downto 0);
	signal P_HR_S37 : unsigned(11 downto 0);
	signal P_HR_S38 : unsigned(11 downto 0);
	signal P_HR_S39 : unsigned(11 downto 0);
	signal P_HR_S40 : unsigned(11 downto 0);
	signal P_HR_S41 : unsigned(11 downto 0);
	signal P_HR_S42 : unsigned(11 downto 0);
	signal P_HR_S43 : unsigned(11 downto 0);
	signal P_HR_S44 : unsigned(11 downto 0);
	signal P_HR_S45 : unsigned(11 downto 0);
	signal P_HR_S46 : unsigned(11 downto 0);
	signal P_HR_S47 : unsigned(11 downto 0);
	signal P_HR_S48 : unsigned(11 downto 0);
	signal P_HR_S49 : unsigned(11 downto 0);
	signal P_HR_S50 : unsigned(11 downto 0);
	signal P_HR_S51 : unsigned(11 downto 0);
	signal P_HR_S52 : unsigned(11 downto 0);
	signal P_HR_S53 : unsigned(11 downto 0);
	signal P_HR_S54 : unsigned(11 downto 0);
	signal P_HR_S55 : unsigned(11 downto 0);
	signal P_HR_S56 : unsigned(11 downto 0);
	signal P_HR_S57 : unsigned(11 downto 0);
	signal P_HR_S58 : unsigned(11 downto 0);
	signal P_HR_S59 : unsigned(11 downto 0);
	signal P_HR_S60 : unsigned(11 downto 0);
	signal P_HR_S61 : unsigned(11 downto 0);
	signal P_HR_S62 : unsigned(11 downto 0);
	signal P_HR_S63 : unsigned(11 downto 0);
	signal P_HR_S64 : unsigned(11 downto 0);
	signal P_HR_S65 : unsigned(11 downto 0);
	signal P_HR_S66 : unsigned(11 downto 0);
	signal P_HR_S67 : unsigned(11 downto 0);
	signal P_HR_S68 : unsigned(11 downto 0);
	signal P_HR_S69 : unsigned(11 downto 0);
	signal P_HR_S70 : unsigned(11 downto 0);
	signal P_HR_S71 : unsigned(11 downto 0);
	signal P_HR_S72 : unsigned(11 downto 0);
	signal P_HR_S73 : unsigned(11 downto 0);
	signal P_HR_S74 : unsigned(11 downto 0);
	signal P_HR_S75 : unsigned(11 downto 0);
	signal P_HR_S76 : unsigned(11 downto 0);
	signal P_HR_S77 : unsigned(11 downto 0);
	signal P_HR_S78 : unsigned(11 downto 0);
	signal P_HR_S79 : unsigned(11 downto 0);
	signal P_HR_S80 : unsigned(11 downto 0);
	signal P_HR_S81 : unsigned(11 downto 0);
	signal P_HR_S82 : unsigned(11 downto 0);
	signal P_HR_S83 : unsigned(11 downto 0);
	signal P_HR_S84 : unsigned(11 downto 0);
	signal P_HR_S85 : unsigned(11 downto 0);
	signal P_HR_S86 : unsigned(11 downto 0);
	signal P_HR_S87 : unsigned(11 downto 0);
	signal P_HR_S88 : unsigned(11 downto 0);
	signal P_HR_S89 : unsigned(11 downto 0);
	signal P_HR_S90 : unsigned(11 downto 0);
	signal P_HR_S91 : unsigned(11 downto 0);
	signal P_HR_S92 : unsigned(11 downto 0);
	signal P_HR_S93 : unsigned(11 downto 0);
	signal P_HR_S94 : unsigned(11 downto 0);
	signal P_HR_S95 : unsigned(11 downto 0);
	signal P_HR_S96 : unsigned(11 downto 0);
	signal P_HR_S97 : unsigned(11 downto 0);
	signal P_HR_S98 : unsigned(11 downto 0);
	signal P_HR_S99 : unsigned(11 downto 0);
	signal P_HR_S100 : unsigned(11 downto 0);
	signal P_HR_S101 : unsigned(11 downto 0);
	signal P_HR_S102 : unsigned(11 downto 0);
	signal P_HR_S103 : unsigned(11 downto 0);
	signal P_HR_S104 : unsigned(11 downto 0);
	signal P_HR_S105 : unsigned(11 downto 0);
	signal P_HR_S106 : unsigned(11 downto 0);
	signal P_HR_S107 : unsigned(11 downto 0);
	signal P_HR_S108 : unsigned(11 downto 0);
	signal P_HR_S109 : unsigned(11 downto 0);
	signal P_HR_S110 : unsigned(11 downto 0);
	signal P_HR_S111 : unsigned(11 downto 0);
	signal P_HR_S112 : unsigned(11 downto 0);
	signal P_HR_S113 : unsigned(11 downto 0);
	signal P_HR_S114 : unsigned(11 downto 0);
	signal P_HR_S115 : unsigned(11 downto 0);
	signal P_HR_S116 : unsigned(11 downto 0);
	signal P_HR_S117 : unsigned(11 downto 0);
	signal P_HR_S118 : unsigned(11 downto 0);
	signal P_HR_S119 : unsigned(11 downto 0);
	signal P_HR_S120 : unsigned(11 downto 0);
	signal P_HR_S121 : unsigned(11 downto 0);
	signal P_HR_S122 : unsigned(11 downto 0);
	signal P_HR_S123 : unsigned(11 downto 0);
	signal P_HR_S124 : unsigned(11 downto 0);
	signal P_HR_S125 : unsigned(11 downto 0);
	signal P_HR_S126 : unsigned(11 downto 0);
	signal P_HR_S127 : unsigned(11 downto 0);
	signal P_HR_S128 : unsigned(11 downto 0);
	signal P_HR_S129 : unsigned(11 downto 0);
	signal P_HR_S130 : unsigned(11 downto 0);
	signal P_HR_S131 : unsigned(11 downto 0);
	signal P_HR_S132 : unsigned(11 downto 0);
	signal P_HR_S133 : unsigned(11 downto 0);
	signal P_HR_S134 : unsigned(11 downto 0);
	signal P_HR_S135 : unsigned(11 downto 0);
	signal P_HR_S136 : unsigned(11 downto 0);
	signal P_HR_S137 : unsigned(11 downto 0);
	signal P_HR_S138 : unsigned(11 downto 0);
	signal P_HR_S139 : unsigned(11 downto 0);
	signal P_HR_S140 : unsigned(11 downto 0);
	signal P_HR_S141 : unsigned(11 downto 0);
	signal P_HR_S142 : unsigned(11 downto 0);
	signal P_HR_S143 : unsigned(11 downto 0);
	signal P_HR_S144 : unsigned(11 downto 0);
	signal P_HR_S145 : unsigned(11 downto 0);
	signal P_HR_S146 : unsigned(11 downto 0);
	signal P_HR_S147 : unsigned(11 downto 0);
	signal P_HR_S148 : unsigned(11 downto 0);
	signal P_HR_S149 : unsigned(11 downto 0);
	signal P_HR_S150 : unsigned(11 downto 0);
	signal P_HR_S151 : unsigned(11 downto 0);
	signal P_HR_S152 : unsigned(11 downto 0);
	signal P_HR_S153 : unsigned(11 downto 0);
	signal P_HR_S154 : unsigned(11 downto 0);
	signal P_HR_S155 : unsigned(11 downto 0);
	signal P_HR_S156 : unsigned(11 downto 0);
	signal P_HR_S157 : unsigned(11 downto 0);
	signal P_HR_S158 : unsigned(11 downto 0);
	signal P_HR_S159 : unsigned(11 downto 0);
	signal P_HR_S160 : unsigned(11 downto 0);
	signal P_HR_S161 : unsigned(11 downto 0);
	signal P_HR_S162 : unsigned(11 downto 0);
	signal P_HR_S163 : unsigned(11 downto 0);
	signal P_HR_S164 : unsigned(11 downto 0);
	signal P_HR_S165 : unsigned(11 downto 0);
	signal P_HR_S166 : unsigned(11 downto 0);
	signal P_HR_S167 : unsigned(11 downto 0);
	signal P_HR_S168 : unsigned(11 downto 0);
	signal P_HR_S169 : unsigned(11 downto 0);
	signal P_HR_S170 : unsigned(11 downto 0);
	signal P_HR_S171 : unsigned(11 downto 0);
	signal P_HR_S172 : unsigned(11 downto 0);
	signal P_HR_S173 : unsigned(11 downto 0);
	signal P_HR_S174 : unsigned(11 downto 0);
	signal P_HR_S175 : unsigned(11 downto 0);
	signal P_HR_S176 : unsigned(11 downto 0);
	signal P_HR_S177 : unsigned(11 downto 0);
	signal P_HR_S178 : unsigned(11 downto 0);
	signal P_HR_S179 : unsigned(11 downto 0);
	signal P_HR_S180 : unsigned(11 downto 0);
	signal P_HR_S181 : unsigned(11 downto 0);
	signal P_HR_S182 : unsigned(11 downto 0);
	signal P_HR_S183 : unsigned(11 downto 0);
	signal P_HR_S184 : unsigned(11 downto 0);
	signal P_HR_S185 : unsigned(11 downto 0);
	signal P_HR_S186 : unsigned(11 downto 0);
	signal P_HR_S187 : unsigned(11 downto 0);
	signal P_HR_S188 : unsigned(11 downto 0);
	signal P_HR_S189 : unsigned(11 downto 0);
	signal P_HR_S190 : unsigned(11 downto 0);
	signal P_HR_S191 : unsigned(11 downto 0);
	signal P_HR_S192 : unsigned(11 downto 0);
	signal P_HR_S193 : unsigned(11 downto 0);
	signal P_HR_S194 : unsigned(11 downto 0);
	signal P_HR_S195 : unsigned(11 downto 0);
	signal P_HR_S196 : unsigned(11 downto 0);
	signal P_HR_S197 : unsigned(11 downto 0);
	signal P_HR_S198 : unsigned(11 downto 0);
	signal P_HR_S199 : unsigned(11 downto 0);
	signal P_HR_S200 : unsigned(11 downto 0);
	signal P_HR_S201 : unsigned(11 downto 0);
	signal P_HR_S202 : unsigned(11 downto 0);
	signal P_HR_S203 : unsigned(11 downto 0);
	signal P_HR_S204 : unsigned(11 downto 0);
	signal P_HR_S205 : unsigned(11 downto 0);
	signal P_HR_S206 : unsigned(11 downto 0);
	signal P_HR_S207 : unsigned(11 downto 0);
	signal P_HR_S208 : unsigned(11 downto 0);
	signal P_HR_S209 : unsigned(11 downto 0);
	signal P_HR_S210 : unsigned(11 downto 0);
	signal P_HR_S211 : unsigned(11 downto 0);
	signal P_HR_S212 : unsigned(11 downto 0);
	signal P_HR_S213 : unsigned(11 downto 0);
	signal P_HR_S214 : unsigned(11 downto 0);
	signal P_HR_S215 : unsigned(11 downto 0);
	signal P_HR_S216 : unsigned(11 downto 0);
	signal P_HR_S217 : unsigned(11 downto 0);
	signal P_HR_S218 : unsigned(11 downto 0);
	signal P_HR_S219 : unsigned(11 downto 0);
	signal P_HR_S220 : unsigned(11 downto 0);
	signal P_HR_S221 : unsigned(11 downto 0);
	signal P_HR_S222 : unsigned(11 downto 0);
	signal P_HR_S223 : unsigned(11 downto 0);
	signal P_HR_S224 : unsigned(11 downto 0);
	signal P_HR_S225 : unsigned(11 downto 0);
	signal P_HR_S226 : unsigned(11 downto 0);
	signal P_HR_S227 : unsigned(11 downto 0);
	signal P_HR_S228 : unsigned(11 downto 0);
	signal P_HR_S229 : unsigned(11 downto 0);
	signal P_HR_S230 : unsigned(11 downto 0);
	signal P_HR_S231 : unsigned(11 downto 0);
	signal P_HR_S232 : unsigned(11 downto 0);
	signal P_HR_S233 : unsigned(11 downto 0);
	signal P_HR_S234 : unsigned(11 downto 0);
	signal P_HR_S235 : unsigned(11 downto 0);
	signal P_HR_S236 : unsigned(11 downto 0);
	signal P_HR_S237 : unsigned(11 downto 0);
	signal P_HR_S238 : unsigned(11 downto 0);
	signal P_HR_S239 : unsigned(11 downto 0);
	signal P_HR_S240 : unsigned(11 downto 0);
	signal P_HR_S241 : unsigned(11 downto 0);
	signal P_HR_S242 : unsigned(11 downto 0);
	signal P_HR_S243 : unsigned(11 downto 0);
	signal P_HR_S244 : unsigned(11 downto 0);
	signal P_HR_S245 : unsigned(11 downto 0);
	signal P_HR_S246 : unsigned(11 downto 0);
	signal P_HR_S247 : unsigned(11 downto 0);
	signal P_HR_S248 : unsigned(11 downto 0);
	signal P_HR_S249 : unsigned(11 downto 0);
	signal P_HR_S250 : unsigned(11 downto 0);
	signal P_HR_S251 : unsigned(11 downto 0);
	signal P_HR_S252 : unsigned(11 downto 0);
	signal P_HR_S253 : unsigned(11 downto 0);
	signal P_HR_S254 : unsigned(11 downto 0);
	signal P_HR_S255 : unsigned(11 downto 0);
	signal P_HR_S256 : unsigned(11 downto 0);
	signal P_HR_S257 : unsigned(11 downto 0);
	signal P_HR_S258 : unsigned(11 downto 0);
	signal P_HR_S259 : unsigned(11 downto 0);
	signal P_HR_S260 : unsigned(11 downto 0);
	signal P_HR_S261 : unsigned(11 downto 0);
	signal P_HR_S262 : unsigned(11 downto 0);
	signal P_HR_S263 : unsigned(11 downto 0);
	signal P_HR_S264 : unsigned(11 downto 0);
	signal P_HR_S265 : unsigned(11 downto 0);
	signal P_HR_S266 : unsigned(11 downto 0);
	signal P_HR_S267 : unsigned(11 downto 0);
	signal P_HR_S268 : unsigned(11 downto 0);
	signal P_HR_S269 : unsigned(11 downto 0);
	signal P_HR_S270 : unsigned(11 downto 0);
	signal P_HR_S271 : unsigned(11 downto 0);
	signal P_HR_S272 : unsigned(11 downto 0);
	signal P_HR_S273 : unsigned(11 downto 0);
	signal P_HR_S274 : unsigned(11 downto 0);
	signal P_HR_S275 : unsigned(11 downto 0);
	signal P_HR_S276 : unsigned(11 downto 0);
	signal P_HR_S277 : unsigned(11 downto 0);
	signal P_HR_S278 : unsigned(11 downto 0);
	signal P_HR_S279 : unsigned(11 downto 0);
	signal P_HR_S280 : unsigned(11 downto 0);
	signal P_HR_S281 : unsigned(11 downto 0);
	signal P_HR_S282 : unsigned(11 downto 0);
	signal P_HR_S283 : unsigned(11 downto 0);
	signal P_HR_S284 : unsigned(11 downto 0);
	signal P_HR_S285 : unsigned(11 downto 0);
	signal P_HR_S286 : unsigned(11 downto 0);
	signal P_HR_S287 : unsigned(11 downto 0);
	signal P_HR_S288 : unsigned(11 downto 0);
	signal P_HR_S289 : unsigned(11 downto 0);
	signal P_HR_S290 : unsigned(11 downto 0);
	signal P_HR_S291 : unsigned(11 downto 0);
	signal P_HR_S292 : unsigned(11 downto 0);
	signal P_HR_S293 : unsigned(11 downto 0);
	signal P_HR_S294 : unsigned(11 downto 0);
	signal P_HR_S295 : unsigned(11 downto 0);
	signal P_HR_S296 : unsigned(11 downto 0);
	signal P_HR_S297 : unsigned(11 downto 0);
	signal P_HR_S298 : unsigned(11 downto 0);
	signal P_HR_S299 : unsigned(11 downto 0);
	signal P_HR_S300 : unsigned(11 downto 0);
	signal P_HR_S301 : unsigned(11 downto 0);
	signal P_HR_S302 : unsigned(11 downto 0);
	signal P_HR_S303 : unsigned(11 downto 0);
	signal P_HR_S304 : unsigned(11 downto 0);
	signal P_HR_S305 : unsigned(11 downto 0);
	signal P_HR_S306 : unsigned(11 downto 0);
	signal P_HR_S307 : unsigned(11 downto 0);
	signal P_HR_S308 : unsigned(11 downto 0);
	signal P_HR_S309 : unsigned(11 downto 0);
	signal P_HR_S310 : unsigned(11 downto 0);
	signal P_HR_S311 : unsigned(11 downto 0);
	signal P_HR_S312 : unsigned(11 downto 0);
	signal P_HR_S313 : unsigned(11 downto 0);
	signal P_HR_S314 : unsigned(11 downto 0);
	signal P_HR_S315 : unsigned(11 downto 0);
	signal P_HR_S316 : unsigned(11 downto 0);
	signal P_HR_S317 : unsigned(11 downto 0);
	signal P_HR_S318 : unsigned(11 downto 0);
	signal P_HR_S319 : unsigned(11 downto 0);
	signal P_HR_S320 : unsigned(11 downto 0);
	signal P_HR_S321 : unsigned(11 downto 0);
	signal P_HR_S322 : unsigned(11 downto 0);
	signal P_HR_S323 : unsigned(11 downto 0);
	signal P_HR_S324 : unsigned(11 downto 0);
	signal P_HR_S325 : unsigned(11 downto 0);
	signal P_HR_S326 : unsigned(11 downto 0);
	signal P_HR_S327 : unsigned(11 downto 0);
	signal P_HR_S328 : unsigned(11 downto 0);
	signal P_HR_S329 : unsigned(11 downto 0);
	signal P_HR_S330 : unsigned(11 downto 0);
	signal P_HR_S331 : unsigned(11 downto 0);
	signal P_HR_S332 : unsigned(11 downto 0);
	signal P_HR_S333 : unsigned(11 downto 0);
	signal P_HR_S334 : unsigned(11 downto 0);
	signal P_HR_S335 : unsigned(11 downto 0);
	signal P_HR_S336 : unsigned(11 downto 0);
	signal P_HR_S337 : unsigned(11 downto 0);
	signal P_HR_S338 : unsigned(11 downto 0);
	signal P_HR_S339 : unsigned(11 downto 0);
	signal P_HR_S340 : unsigned(11 downto 0);
	signal P_HR_S341 : unsigned(11 downto 0);
	signal P_HR_S342 : unsigned(11 downto 0);
	signal P_HR_S343 : unsigned(11 downto 0);
	signal P_HR_S344 : unsigned(11 downto 0);
	signal P_HR_S345 : unsigned(11 downto 0);
	signal P_HR_S346 : unsigned(11 downto 0);
	signal P_HR_S347 : unsigned(11 downto 0);
	signal P_HR_S348 : unsigned(11 downto 0);
	signal P_HR_S349 : unsigned(11 downto 0);
	signal P_HR_S350 : unsigned(11 downto 0);
	signal P_HR_S351 : unsigned(11 downto 0);
	signal P_HR_S352 : unsigned(11 downto 0);
	signal P_HR_S353 : unsigned(11 downto 0);
	signal P_HR_S354 : unsigned(11 downto 0);
	signal P_HR_S355 : unsigned(11 downto 0);
	signal P_HR_S356 : unsigned(11 downto 0);
	signal P_HR_S357 : unsigned(11 downto 0);
	signal P_HR_S358 : unsigned(11 downto 0);
	signal P_HR_S359 : unsigned(11 downto 0);
	signal P_HR_S360 : unsigned(11 downto 0);
	signal P_HR_S361 : unsigned(11 downto 0);
	signal P_HR_S362 : unsigned(11 downto 0);
	signal P_HR_S363 : unsigned(11 downto 0);
	signal P_HR_S364 : unsigned(11 downto 0);
	signal P_HR_S365 : unsigned(11 downto 0);
	signal P_HR_S366 : unsigned(11 downto 0);
	signal P_HR_S367 : unsigned(11 downto 0);
	signal P_HR_S368 : unsigned(11 downto 0);
	signal P_HR_S369 : unsigned(11 downto 0);
	signal P_HR_S370 : unsigned(11 downto 0);
	signal P_HR_S371 : unsigned(11 downto 0);
	signal P_HR_S372 : unsigned(11 downto 0);
	signal P_HR_S373 : unsigned(11 downto 0);
	signal P_HR_S374 : unsigned(11 downto 0);
	signal P_HR_S375 : unsigned(11 downto 0);
	signal P_HR_S376 : unsigned(11 downto 0);
	signal P_HR_S377 : unsigned(11 downto 0);
	signal P_HR_S378 : unsigned(11 downto 0);
	signal P_HR_S379 : unsigned(11 downto 0);
	signal P_HR_S380 : unsigned(11 downto 0);
	signal P_HR_S381 : unsigned(11 downto 0);
	signal P_HR_S382 : unsigned(11 downto 0);
	signal P_HR_S383 : unsigned(11 downto 0);
	signal P_HR_S384 : unsigned(11 downto 0);
	signal P_HR_S385 : unsigned(11 downto 0);
	signal P_HR_S386 : unsigned(11 downto 0);
	signal P_HR_S387 : unsigned(11 downto 0);
	signal P_HR_S388 : unsigned(11 downto 0);
	signal P_HR_S389 : unsigned(11 downto 0);
	signal P_HR_S390 : unsigned(11 downto 0);
	signal P_HR_S391 : unsigned(11 downto 0);
	signal P_HR_S392 : unsigned(11 downto 0);
	signal P_HR_S393 : unsigned(11 downto 0);
	signal P_HR_S394 : unsigned(11 downto 0);
	signal P_HR_S395 : unsigned(11 downto 0);
	signal P_HR_S396 : unsigned(11 downto 0);
	signal P_HR_S397 : unsigned(11 downto 0);
	signal P_HR_S398 : unsigned(11 downto 0);
	signal P_HR_S399 : unsigned(11 downto 0);
	signal P_HR_S400 : unsigned(11 downto 0);
	signal P_HR_S401 : unsigned(11 downto 0);
	signal P_HR_S402 : unsigned(11 downto 0);
	signal P_HR_S403 : unsigned(11 downto 0);
	signal P_HR_S404 : unsigned(11 downto 0);
	signal P_HR_S405 : unsigned(11 downto 0);
	signal P_HR_S406 : unsigned(11 downto 0);
	signal P_HR_S407 : unsigned(11 downto 0);
	signal P_HR_S408 : unsigned(11 downto 0);
	signal P_HR_S409 : unsigned(11 downto 0);
	signal P_HR_S410 : unsigned(11 downto 0);
	signal P_HR_S411 : unsigned(11 downto 0);
	signal P_HR_S412 : unsigned(11 downto 0);
	signal P_HR_S413 : unsigned(11 downto 0);
	signal P_HR_S414 : unsigned(11 downto 0);
	signal P_HR_S415 : unsigned(11 downto 0);
	signal P_HR_S416 : unsigned(11 downto 0);
	signal P_HR_S417 : unsigned(11 downto 0);
	signal P_HR_S418 : unsigned(11 downto 0);
	signal P_HR_S419 : unsigned(11 downto 0);
	signal P_HR_S420 : unsigned(11 downto 0);
	signal P_HR_S421 : unsigned(11 downto 0);
	signal P_HR_S422 : unsigned(11 downto 0);
	signal P_HR_S423 : unsigned(11 downto 0);
	signal P_HR_S424 : unsigned(11 downto 0);
	signal P_HR_S425 : unsigned(11 downto 0);
	signal P_HR_S426 : unsigned(11 downto 0);
	signal P_HR_S427 : unsigned(11 downto 0);
	signal P_HR_S428 : unsigned(11 downto 0);
	signal P_HR_S429 : unsigned(11 downto 0);
	signal P_HR_S430 : unsigned(11 downto 0);
	signal P_HR_S431 : unsigned(11 downto 0);
	signal P_HR_S432 : unsigned(11 downto 0);
	signal P_HR_S433 : unsigned(11 downto 0);
	signal P_HR_S434 : unsigned(11 downto 0);
	signal P_HR_S435 : unsigned(11 downto 0);
	signal P_HR_S436 : unsigned(11 downto 0);
	signal P_HR_S437 : unsigned(11 downto 0);
	signal P_HR_S438 : unsigned(11 downto 0);
	signal P_HR_S439 : unsigned(11 downto 0);
	signal P_HR_S440 : unsigned(11 downto 0);
	signal P_HR_S441 : unsigned(11 downto 0);
	signal P_HR_S442 : unsigned(11 downto 0);
	signal P_HR_S443 : unsigned(11 downto 0);
	signal P_HR_S444 : unsigned(11 downto 0);
	signal P_HR_S445 : unsigned(11 downto 0);
	signal P_HR_S446 : unsigned(11 downto 0);
	signal P_HR_S447 : unsigned(11 downto 0);
	signal P_HR_S448 : unsigned(11 downto 0);
	signal P_HR_S449 : unsigned(11 downto 0);
	signal P_HR_S450 : unsigned(11 downto 0);
	signal P_HR_S451 : unsigned(11 downto 0);
	signal P_HR_S452 : unsigned(11 downto 0);
	signal P_HR_S453 : unsigned(11 downto 0);
	signal P_HR_S454 : unsigned(11 downto 0);
	signal P_HR_S455 : unsigned(11 downto 0);
	signal P_HR_S456 : unsigned(11 downto 0);
	signal P_HR_S457 : unsigned(11 downto 0);
	signal P_HR_S458 : unsigned(11 downto 0);
	signal P_HR_S459 : unsigned(11 downto 0);
	signal P_HR_S460 : unsigned(11 downto 0);
	signal P_HR_S461 : unsigned(11 downto 0);
	signal P_HR_S462 : unsigned(11 downto 0);
	signal P_HR_S463 : unsigned(11 downto 0);
	signal P_HR_S464 : unsigned(11 downto 0);
	signal P_HR_S465 : unsigned(11 downto 0);
	signal P_HR_S466 : unsigned(11 downto 0);
	signal P_HR_S467 : unsigned(11 downto 0);
	signal P_HR_S468 : unsigned(11 downto 0);
	signal P_HR_S469 : unsigned(11 downto 0);
	signal P_HR_S470 : unsigned(11 downto 0);
	signal P_HR_S471 : unsigned(11 downto 0);
	signal P_HR_S472 : unsigned(11 downto 0);
	signal P_HR_S473 : unsigned(11 downto 0);
	signal P_HR_S474 : unsigned(11 downto 0);
	signal P_HR_S475 : unsigned(11 downto 0);
	signal P_HR_S476 : unsigned(11 downto 0);
	signal P_HR_S477 : unsigned(11 downto 0);
	signal P_HR_S478 : unsigned(11 downto 0);
	signal P_HR_S479 : unsigned(11 downto 0);
	signal P_HR_S480 : unsigned(11 downto 0);
	signal P_HR_S481 : unsigned(11 downto 0);
	signal P_HR_S482 : unsigned(11 downto 0);
	signal P_HR_S483 : unsigned(11 downto 0);
	signal P_HR_S484 : unsigned(11 downto 0);
	signal P_HR_S485 : unsigned(11 downto 0);
	signal P_HR_S486 : unsigned(11 downto 0);
	signal P_HR_S487 : unsigned(11 downto 0);
	signal P_HR_S488 : unsigned(11 downto 0);
	signal P_HR_S489 : unsigned(11 downto 0);
	signal P_HR_S490 : unsigned(11 downto 0);
	signal P_HR_S491 : unsigned(11 downto 0);
	signal P_HR_S492 : unsigned(11 downto 0);
	signal P_HR_S493 : unsigned(11 downto 0);
	signal P_HR_S494 : unsigned(11 downto 0);
	signal P_HR_S495 : unsigned(11 downto 0);
	signal P_HR_S496 : unsigned(11 downto 0);
	signal P_HR_S497 : unsigned(11 downto 0);
	signal P_HR_S498 : unsigned(11 downto 0);
	signal P_HR_S499 : unsigned(11 downto 0);
	signal P_HR_S500 : unsigned(11 downto 0);
	signal P_HR_S501 : unsigned(11 downto 0);
	signal P_HR_S502 : unsigned(11 downto 0);
	signal P_HR_S503 : unsigned(11 downto 0);
	signal P_HR_S504 : unsigned(11 downto 0);
	signal P_HR_S505 : unsigned(11 downto 0);
	signal P_HR_S506 : unsigned(11 downto 0);
	signal P_HR_S507 : unsigned(11 downto 0);
	signal P_HR_S508 : unsigned(11 downto 0);
	signal P_HR_S509 : unsigned(11 downto 0);
	signal P_HR_S510 : unsigned(11 downto 0);
	signal P_HR_S511 : unsigned(11 downto 0);
	signal P_HR_S512 : unsigned(11 downto 0);
	signal P_HR_S513 : unsigned(11 downto 0);
	signal P_HR_S514 : unsigned(11 downto 0);
	signal P_HR_S515 : unsigned(11 downto 0);
	signal P_HR_S516 : unsigned(11 downto 0);
	signal P_HR_S517 : unsigned(11 downto 0);
	signal P_HR_S518 : unsigned(11 downto 0);
	signal P_HR_S519 : unsigned(11 downto 0);
	signal P_HR_S520 : unsigned(11 downto 0);
	signal P_HR_S521 : unsigned(11 downto 0);
	signal P_HR_S522 : unsigned(11 downto 0);
	signal P_HR_S523 : unsigned(11 downto 0);
	signal P_HR_S524 : unsigned(11 downto 0);
	signal P_HR_S525 : unsigned(11 downto 0);
	signal P_HR_S526 : unsigned(11 downto 0);
	signal P_HR_S527 : unsigned(11 downto 0);
	signal P_HR_S528 : unsigned(11 downto 0);
	signal P_HR_S529 : unsigned(11 downto 0);
	signal P_HR_S530 : unsigned(11 downto 0);
	signal P_HR_S531 : unsigned(11 downto 0);
	signal P_HR_S532 : unsigned(11 downto 0);
	signal P_HR_S533 : unsigned(11 downto 0);
	signal P_HR_S534 : unsigned(11 downto 0);
	signal P_HR_S535 : unsigned(11 downto 0);
	signal P_HR_S536 : unsigned(11 downto 0);
	signal P_HR_S537 : unsigned(11 downto 0);
	signal P_HR_S538 : unsigned(11 downto 0);
	signal P_HR_S539 : unsigned(11 downto 0);
	signal P_HR_S540 : unsigned(11 downto 0);
	signal P_HR_S541 : unsigned(11 downto 0);
	signal P_HR_S542 : unsigned(11 downto 0);
	signal P_HR_S543 : unsigned(11 downto 0);
	signal P_HR_S544 : unsigned(11 downto 0);
	signal P_HR_S545 : unsigned(11 downto 0);
	signal P_HR_S546 : unsigned(11 downto 0);
	signal P_HR_S547 : unsigned(11 downto 0);
	signal P_HR_S548 : unsigned(11 downto 0);
	signal P_HR_S549 : unsigned(11 downto 0);
	signal P_HR_S550 : unsigned(11 downto 0);
	signal P_HR_S551 : unsigned(11 downto 0);
	signal P_HR_S552 : unsigned(11 downto 0);
	signal P_HR_S553 : unsigned(11 downto 0);
	signal P_HR_S554 : unsigned(11 downto 0);
	signal P_HR_S555 : unsigned(11 downto 0);
	signal P_HR_S556 : unsigned(11 downto 0);
	signal P_HR_S557 : unsigned(11 downto 0);
	signal P_HR_S558 : unsigned(11 downto 0);
	signal P_HR_S559 : unsigned(11 downto 0);
	signal P_HR_S560 : unsigned(11 downto 0);
	signal P_HR_S561 : unsigned(11 downto 0);
	signal P_HR_S562 : unsigned(11 downto 0);
	signal P_HR_S563 : unsigned(11 downto 0);
	signal P_HR_S564 : unsigned(11 downto 0);
	signal P_HR_S565 : unsigned(11 downto 0);
	signal P_HR_S566 : unsigned(11 downto 0);
	signal P_HR_S567 : unsigned(11 downto 0);
	signal P_HR_S568 : unsigned(11 downto 0);
	signal P_HR_S569 : unsigned(11 downto 0);
	signal P_HR_S570 : unsigned(11 downto 0);
	signal P_HR_S571 : unsigned(11 downto 0);
	signal P_HR_S572 : unsigned(11 downto 0);
	signal P_HR_S573 : unsigned(11 downto 0);
	signal P_HR_S574 : unsigned(11 downto 0);
	signal P_HR_S575 : unsigned(11 downto 0);
	signal P_HR_S576 : unsigned(11 downto 0);
	signal P_HR_S577 : unsigned(11 downto 0);
	signal P_HR_S578 : unsigned(11 downto 0);
	signal P_HR_S579 : unsigned(11 downto 0);
	signal P_HR_S580 : unsigned(11 downto 0);
	signal P_HR_S581 : unsigned(11 downto 0);
	signal P_HR_S582 : unsigned(11 downto 0);
	signal P_HR_S583 : unsigned(11 downto 0);
	signal P_HR_S584 : unsigned(11 downto 0);
	signal P_HR_S585 : unsigned(11 downto 0);
	signal P_HR_S586 : unsigned(11 downto 0);
	signal P_HR_S587 : unsigned(11 downto 0);
	signal P_HR_S588 : unsigned(11 downto 0);
	signal P_HR_S589 : unsigned(11 downto 0);
	signal P_HR_S590 : unsigned(11 downto 0);
	signal P_HR_S591 : unsigned(11 downto 0);
	signal P_HR_S592 : unsigned(11 downto 0);
	signal P_HR_S593 : unsigned(11 downto 0);
	signal P_HR_S594 : unsigned(11 downto 0);
	signal P_HR_S595 : unsigned(11 downto 0);
	signal P_HR_S596 : unsigned(11 downto 0);
	signal P_HR_S597 : unsigned(11 downto 0);
	signal P_HR_S598 : unsigned(11 downto 0);
	signal P_HR_S599 : unsigned(11 downto 0);
	signal P_HR_S600 : unsigned(11 downto 0);
	signal P_HR_S601 : unsigned(11 downto 0);
	signal P_HR_S602 : unsigned(11 downto 0);
	signal P_HR_S603 : unsigned(11 downto 0);
	signal P_HR_S604 : unsigned(11 downto 0);
	signal P_HR_S605 : unsigned(11 downto 0);
	signal P_HR_S606 : unsigned(11 downto 0);
	signal P_HR_S607 : unsigned(11 downto 0);
	signal P_HR_S608 : unsigned(11 downto 0);
	signal P_HR_S609 : unsigned(11 downto 0);
	signal P_HR_S610 : unsigned(11 downto 0);
	signal P_HR_S611 : unsigned(11 downto 0);
	signal P_HR_S612 : unsigned(11 downto 0);
	signal P_HR_S613 : unsigned(11 downto 0);
	signal P_HR_S614 : unsigned(11 downto 0);
	signal P_HR_S615 : unsigned(11 downto 0);
	signal P_HR_S616 : unsigned(11 downto 0);
	signal P_HR_S617 : unsigned(11 downto 0);
	signal P_HR_S618 : unsigned(11 downto 0);
	signal P_HR_S619 : unsigned(11 downto 0);
	signal P_HR_S620 : unsigned(11 downto 0);
	signal P_HR_S621 : unsigned(11 downto 0);
	signal P_HR_S622 : unsigned(11 downto 0);
	signal P_HR_S623 : unsigned(11 downto 0);
	signal P_HR_S624 : unsigned(11 downto 0);
	
	
    signal P_TEMP_NS1 : unsigned(11 downto 0);
    signal P_TEMP_NS2 : unsigned(11 downto 0);
    signal P_TEMP_NS3 : unsigned(11 downto 0);
    signal P_TEMP_NS4 : unsigned(11 downto 0);
    signal P_TEMP_NS5 : unsigned(11 downto 0);
    signal P_TEMP_NS6 : unsigned(11 downto 0);
    signal P_TEMP_NS7 : unsigned(11 downto 0);
    signal P_TEMP_NS8 : unsigned(11 downto 0);
    signal P_TEMP_NS9 : unsigned(11 downto 0);
    signal P_TEMP_NS10 : unsigned(11 downto 0);
    signal P_TEMP_NS11 : unsigned(11 downto 0);
    signal P_TEMP_NS12 : unsigned(11 downto 0);
    signal P_TEMP_NS13 : unsigned(11 downto 0);
    signal P_TEMP_NS14 : unsigned(11 downto 0);
    signal P_TEMP_NS15 : unsigned(11 downto 0);
    signal P_TEMP_NS16 : unsigned(11 downto 0);
    signal P_TEMP_NS17 : unsigned(11 downto 0);
    signal P_TEMP_NS18 : unsigned(11 downto 0);
    signal P_TEMP_NS19 : unsigned(11 downto 0);
    signal P_TEMP_NS20 : unsigned(11 downto 0);
    signal P_TEMP_NS21 : unsigned(11 downto 0);
    signal P_TEMP_NS22 : unsigned(11 downto 0);
    signal P_TEMP_NS23 : unsigned(11 downto 0);
    signal P_TEMP_NS24 : unsigned(11 downto 0);
    signal P_TEMP_NS25 : unsigned(11 downto 0);
    signal P_TEMP_NS26 : unsigned(11 downto 0);
    signal P_TEMP_NS27 : unsigned(11 downto 0);
    signal P_TEMP_NS28 : unsigned(11 downto 0);
    signal P_TEMP_NS29 : unsigned(11 downto 0);
    signal P_TEMP_NS30 : unsigned(11 downto 0);
    signal P_TEMP_NS31 : unsigned(11 downto 0);
    signal P_TEMP_NS32 : unsigned(11 downto 0);
    signal P_TEMP_NS33 : unsigned(11 downto 0);
    signal P_TEMP_NS34 : unsigned(11 downto 0);
    signal P_TEMP_NS35 : unsigned(11 downto 0);
    signal P_TEMP_NS36 : unsigned(11 downto 0);
    signal P_TEMP_NS37 : unsigned(11 downto 0);
    signal P_TEMP_NS38 : unsigned(11 downto 0);
    signal P_TEMP_NS39 : unsigned(11 downto 0);
    signal P_TEMP_NS40 : unsigned(11 downto 0);
    signal P_TEMP_NS41 : unsigned(11 downto 0);
    signal P_TEMP_NS42 : unsigned(11 downto 0);
    signal P_TEMP_NS43 : unsigned(11 downto 0);
    signal P_TEMP_NS44 : unsigned(11 downto 0);
    signal P_TEMP_NS45 : unsigned(11 downto 0);
    signal P_TEMP_NS46 : unsigned(11 downto 0);
    signal P_TEMP_NS47 : unsigned(11 downto 0);
    signal P_TEMP_NS48 : unsigned(11 downto 0);
    signal P_TEMP_NS49 : unsigned(11 downto 0);
    signal P_TEMP_NS50 : unsigned(11 downto 0);
    signal P_TEMP_NS51 : unsigned(11 downto 0);
    signal P_TEMP_NS52 : unsigned(11 downto 0);
    signal P_TEMP_NS53 : unsigned(11 downto 0);
    signal P_TEMP_NS54 : unsigned(11 downto 0);
    signal P_TEMP_NS55 : unsigned(11 downto 0);
    signal P_TEMP_NS56 : unsigned(11 downto 0);
    signal P_TEMP_NS57 : unsigned(11 downto 0);
    signal P_TEMP_NS58 : unsigned(11 downto 0);
    signal P_TEMP_NS59 : unsigned(11 downto 0);
    signal P_TEMP_NS60 : unsigned(11 downto 0);
    signal P_TEMP_NS61 : unsigned(11 downto 0);
    signal P_TEMP_NS62 : unsigned(11 downto 0);
    signal P_TEMP_NS63 : unsigned(11 downto 0);
		
    signal P_HR_NS1 : unsigned(11 downto 0);
    signal P_HR_NS2 : unsigned(11 downto 0);
    signal P_HR_NS3 : unsigned(11 downto 0);
    signal P_HR_NS4 : unsigned(11 downto 0);
    signal P_HR_NS5 : unsigned(11 downto 0);
    signal P_HR_NS6 : unsigned(11 downto 0);
    signal P_HR_NS7 : unsigned(11 downto 0);
    signal P_HR_NS8 : unsigned(11 downto 0);
    signal P_HR_NS9 : unsigned(11 downto 0);
    signal P_HR_NS10 : unsigned(11 downto 0);
    signal P_HR_NS11 : unsigned(11 downto 0);
    signal P_HR_NS12 : unsigned(11 downto 0);
    signal P_HR_NS13 : unsigned(11 downto 0);
    signal P_HR_NS14 : unsigned(11 downto 0);
    signal P_HR_NS15 : unsigned(11 downto 0);
    signal P_HR_NS16 : unsigned(11 downto 0);
    signal P_HR_NS17 : unsigned(11 downto 0);
    signal P_HR_NS18 : unsigned(11 downto 0);
    signal P_HR_NS19 : unsigned(11 downto 0);
    signal P_HR_NS20 : unsigned(11 downto 0);
    signal P_HR_NS21 : unsigned(11 downto 0);
    signal P_HR_NS22 : unsigned(11 downto 0);
    signal P_HR_NS23 : unsigned(11 downto 0);
    signal P_HR_NS24 : unsigned(11 downto 0);
    signal P_HR_NS25 : unsigned(11 downto 0);
    signal P_HR_NS26 : unsigned(11 downto 0);
    signal P_HR_NS27 : unsigned(11 downto 0);
    signal P_HR_NS28 : unsigned(11 downto 0);
    signal P_HR_NS29 : unsigned(11 downto 0);
    signal P_HR_NS30 : unsigned(11 downto 0);
    signal P_HR_NS31 : unsigned(11 downto 0);
    signal P_HR_NS32 : unsigned(11 downto 0);
    signal P_HR_NS33 : unsigned(11 downto 0);
    signal P_HR_NS34 : unsigned(11 downto 0);
    signal P_HR_NS35 : unsigned(11 downto 0);
    signal P_HR_NS36 : unsigned(11 downto 0);
    signal P_HR_NS37 : unsigned(11 downto 0);
    signal P_HR_NS38 : unsigned(11 downto 0);
    signal P_HR_NS39 : unsigned(11 downto 0);
    signal P_HR_NS40 : unsigned(11 downto 0);
    signal P_HR_NS41 : unsigned(11 downto 0);
    signal P_HR_NS42 : unsigned(11 downto 0);
    signal P_HR_NS43 : unsigned(11 downto 0);
    signal P_HR_NS44 : unsigned(11 downto 0);
    signal P_HR_NS45 : unsigned(11 downto 0);
    signal P_HR_NS46 : unsigned(11 downto 0);
    signal P_HR_NS47 : unsigned(11 downto 0);
    signal P_HR_NS48 : unsigned(11 downto 0);
    signal P_HR_NS49 : unsigned(11 downto 0);
    signal P_HR_NS50 : unsigned(11 downto 0);
    signal P_HR_NS51 : unsigned(11 downto 0);
    signal P_HR_NS52 : unsigned(11 downto 0);
    signal P_HR_NS53 : unsigned(11 downto 0);
    signal P_HR_NS54 : unsigned(11 downto 0);
    signal P_HR_NS55 : unsigned(11 downto 0);
    signal P_HR_NS56 : unsigned(11 downto 0);
    signal P_HR_NS57 : unsigned(11 downto 0);
    signal P_HR_NS58 : unsigned(11 downto 0);
    signal P_HR_NS59 : unsigned(11 downto 0);
    signal P_HR_NS60 : unsigned(11 downto 0);
    signal P_HR_NS61 : unsigned(11 downto 0);
    signal P_HR_NS62 : unsigned(11 downto 0);
    signal P_HR_NS63 : unsigned(11 downto 0);
    signal P_HR_NS64 : unsigned(11 downto 0);
    signal P_HR_NS65 : unsigned(11 downto 0);
    signal P_HR_NS66 : unsigned(11 downto 0);
    signal P_HR_NS67 : unsigned(11 downto 0);
    signal P_HR_NS68 : unsigned(11 downto 0);
    signal P_HR_NS69 : unsigned(11 downto 0);
    signal P_HR_NS70 : unsigned(11 downto 0);
    signal P_HR_NS71 : unsigned(11 downto 0);
    signal P_HR_NS72 : unsigned(11 downto 0);
    signal P_HR_NS73 : unsigned(11 downto 0);
    signal P_HR_NS74 : unsigned(11 downto 0);
    signal P_HR_NS75 : unsigned(11 downto 0);
    signal P_HR_NS76 : unsigned(11 downto 0);
    signal P_HR_NS77 : unsigned(11 downto 0);
    signal P_HR_NS78 : unsigned(11 downto 0);
    signal P_HR_NS79 : unsigned(11 downto 0);
    signal P_HR_NS80 : unsigned(11 downto 0);
    signal P_HR_NS81 : unsigned(11 downto 0);
    signal P_HR_NS82 : unsigned(11 downto 0);
    signal P_HR_NS83 : unsigned(11 downto 0);
    signal P_HR_NS84 : unsigned(11 downto 0);
    signal P_HR_NS85 : unsigned(11 downto 0);
    signal P_HR_NS86 : unsigned(11 downto 0);
    signal P_HR_NS87 : unsigned(11 downto 0);
    signal P_HR_NS88 : unsigned(11 downto 0);
    signal P_HR_NS89 : unsigned(11 downto 0);
    signal P_HR_NS90 : unsigned(11 downto 0);
    signal P_HR_NS91 : unsigned(11 downto 0);
    signal P_HR_NS92 : unsigned(11 downto 0);
    signal P_HR_NS93 : unsigned(11 downto 0);
    signal P_HR_NS94 : unsigned(11 downto 0);
    signal P_HR_NS95 : unsigned(11 downto 0);
    signal P_HR_NS96 : unsigned(11 downto 0);
    signal P_HR_NS97 : unsigned(11 downto 0);
    signal P_HR_NS98 : unsigned(11 downto 0);
    signal P_HR_NS99 : unsigned(11 downto 0);
    signal P_HR_NS100 : unsigned(11 downto 0);
    signal P_HR_NS101 : unsigned(11 downto 0);
    signal P_HR_NS102 : unsigned(11 downto 0);
    signal P_HR_NS103 : unsigned(11 downto 0);
    signal P_HR_NS104 : unsigned(11 downto 0);
    signal P_HR_NS105 : unsigned(11 downto 0);
    signal P_HR_NS106 : unsigned(11 downto 0);
    signal P_HR_NS107 : unsigned(11 downto 0);
    signal P_HR_NS108 : unsigned(11 downto 0);
    signal P_HR_NS109 : unsigned(11 downto 0);
    signal P_HR_NS110 : unsigned(11 downto 0);
    signal P_HR_NS111 : unsigned(11 downto 0);
    signal P_HR_NS112 : unsigned(11 downto 0);
    signal P_HR_NS113 : unsigned(11 downto 0);
    signal P_HR_NS114 : unsigned(11 downto 0);
    signal P_HR_NS115 : unsigned(11 downto 0);
    signal P_HR_NS116 : unsigned(11 downto 0);
    signal P_HR_NS117 : unsigned(11 downto 0);
    signal P_HR_NS118 : unsigned(11 downto 0);
    signal P_HR_NS119 : unsigned(11 downto 0);
    signal P_HR_NS120 : unsigned(11 downto 0);
    signal P_HR_NS121 : unsigned(11 downto 0);
    signal P_HR_NS122 : unsigned(11 downto 0);
    signal P_HR_NS123 : unsigned(11 downto 0);
    signal P_HR_NS124 : unsigned(11 downto 0);
    signal P_HR_NS125 : unsigned(11 downto 0);
    signal P_HR_NS126 : unsigned(11 downto 0);
    signal P_HR_NS127 : unsigned(11 downto 0);
    signal P_HR_NS128 : unsigned(11 downto 0);
    signal P_HR_NS129 : unsigned(11 downto 0);
    signal P_HR_NS130 : unsigned(11 downto 0);
    signal P_HR_NS131 : unsigned(11 downto 0);
    signal P_HR_NS132 : unsigned(11 downto 0);
    signal P_HR_NS133 : unsigned(11 downto 0);
    signal P_HR_NS134 : unsigned(11 downto 0);
    signal P_HR_NS135 : unsigned(11 downto 0);
    signal P_HR_NS136 : unsigned(11 downto 0);
    signal P_HR_NS137 : unsigned(11 downto 0);
    signal P_HR_NS138 : unsigned(11 downto 0);
    signal P_HR_NS139 : unsigned(11 downto 0);
    signal P_HR_NS140 : unsigned(11 downto 0);
    signal P_HR_NS141 : unsigned(11 downto 0);
    signal P_HR_NS142 : unsigned(11 downto 0);
    signal P_HR_NS143 : unsigned(11 downto 0);
    signal P_HR_NS144 : unsigned(11 downto 0);
    signal P_HR_NS145 : unsigned(11 downto 0);
    signal P_HR_NS146 : unsigned(11 downto 0);
    signal P_HR_NS147 : unsigned(11 downto 0);
    signal P_HR_NS148 : unsigned(11 downto 0);
    signal P_HR_NS149 : unsigned(11 downto 0);
    signal P_HR_NS150 : unsigned(11 downto 0);
    signal P_HR_NS151 : unsigned(11 downto 0);
    signal P_HR_NS152 : unsigned(11 downto 0);
    signal P_HR_NS153 : unsigned(11 downto 0);
    signal P_HR_NS154 : unsigned(11 downto 0);
    signal P_HR_NS155 : unsigned(11 downto 0);
    signal P_HR_NS156 : unsigned(11 downto 0);
    signal P_HR_NS157 : unsigned(11 downto 0);
    signal P_HR_NS158 : unsigned(11 downto 0);
    signal P_HR_NS159 : unsigned(11 downto 0);
    signal P_HR_NS160 : unsigned(11 downto 0);
    signal P_HR_NS161 : unsigned(11 downto 0);
    signal P_HR_NS162 : unsigned(11 downto 0);
    signal P_HR_NS163 : unsigned(11 downto 0);
    signal P_HR_NS164 : unsigned(11 downto 0);
    signal P_HR_NS165 : unsigned(11 downto 0);
    signal P_HR_NS166 : unsigned(11 downto 0);
    signal P_HR_NS167 : unsigned(11 downto 0);
    signal P_HR_NS168 : unsigned(11 downto 0);
    signal P_HR_NS169 : unsigned(11 downto 0);
    signal P_HR_NS170 : unsigned(11 downto 0);
    signal P_HR_NS171 : unsigned(11 downto 0);
    signal P_HR_NS172 : unsigned(11 downto 0);
    signal P_HR_NS173 : unsigned(11 downto 0);
    signal P_HR_NS174 : unsigned(11 downto 0);
    signal P_HR_NS175 : unsigned(11 downto 0);
    signal P_HR_NS176 : unsigned(11 downto 0);
    signal P_HR_NS177 : unsigned(11 downto 0);
    signal P_HR_NS178 : unsigned(11 downto 0);
    signal P_HR_NS179 : unsigned(11 downto 0);
    signal P_HR_NS180 : unsigned(11 downto 0);
    signal P_HR_NS181 : unsigned(11 downto 0);
    signal P_HR_NS182 : unsigned(11 downto 0);
    signal P_HR_NS183 : unsigned(11 downto 0);
    signal P_HR_NS184 : unsigned(11 downto 0);
    signal P_HR_NS185 : unsigned(11 downto 0);
    signal P_HR_NS186 : unsigned(11 downto 0);
    signal P_HR_NS187 : unsigned(11 downto 0);
    signal P_HR_NS188 : unsigned(11 downto 0);
    signal P_HR_NS189 : unsigned(11 downto 0);
    signal P_HR_NS190 : unsigned(11 downto 0);
    signal P_HR_NS191 : unsigned(11 downto 0);
    signal P_HR_NS192 : unsigned(11 downto 0);
    signal P_HR_NS193 : unsigned(11 downto 0);
    signal P_HR_NS194 : unsigned(11 downto 0);
    signal P_HR_NS195 : unsigned(11 downto 0);
    signal P_HR_NS196 : unsigned(11 downto 0);
    signal P_HR_NS197 : unsigned(11 downto 0);
    signal P_HR_NS198 : unsigned(11 downto 0);
    signal P_HR_NS199 : unsigned(11 downto 0);
    signal P_HR_NS200 : unsigned(11 downto 0);
    signal P_HR_NS201 : unsigned(11 downto 0);
    signal P_HR_NS202 : unsigned(11 downto 0);
    signal P_HR_NS203 : unsigned(11 downto 0);
    signal P_HR_NS204 : unsigned(11 downto 0);
    signal P_HR_NS205 : unsigned(11 downto 0);
    signal P_HR_NS206 : unsigned(11 downto 0);
    signal P_HR_NS207 : unsigned(11 downto 0);
    signal P_HR_NS208 : unsigned(11 downto 0);
    signal P_HR_NS209 : unsigned(11 downto 0);
    signal P_HR_NS210 : unsigned(11 downto 0);
    signal P_HR_NS211 : unsigned(11 downto 0);
    signal P_HR_NS212 : unsigned(11 downto 0);
    signal P_HR_NS213 : unsigned(11 downto 0);
    signal P_HR_NS214 : unsigned(11 downto 0);
    signal P_HR_NS215 : unsigned(11 downto 0);
    signal P_HR_NS216 : unsigned(11 downto 0);
    signal P_HR_NS217 : unsigned(11 downto 0);
    signal P_HR_NS218 : unsigned(11 downto 0);
    signal P_HR_NS219 : unsigned(11 downto 0);
    signal P_HR_NS220 : unsigned(11 downto 0);
    signal P_HR_NS221 : unsigned(11 downto 0);
    signal P_HR_NS222 : unsigned(11 downto 0);
    signal P_HR_NS223 : unsigned(11 downto 0);
    signal P_HR_NS224 : unsigned(11 downto 0);
    signal P_HR_NS225 : unsigned(11 downto 0);
    signal P_HR_NS226 : unsigned(11 downto 0);
    signal P_HR_NS227 : unsigned(11 downto 0);
    signal P_HR_NS228 : unsigned(11 downto 0);
    signal P_HR_NS229 : unsigned(11 downto 0);
    signal P_HR_NS230 : unsigned(11 downto 0);
    signal P_HR_NS231 : unsigned(11 downto 0);
    signal P_HR_NS232 : unsigned(11 downto 0);
    signal P_HR_NS233 : unsigned(11 downto 0);
    signal P_HR_NS234 : unsigned(11 downto 0);
    signal P_HR_NS235 : unsigned(11 downto 0);
    signal P_HR_NS236 : unsigned(11 downto 0);
    signal P_HR_NS237 : unsigned(11 downto 0);
    signal P_HR_NS238 : unsigned(11 downto 0);
    signal P_HR_NS239 : unsigned(11 downto 0);
    signal P_HR_NS240 : unsigned(11 downto 0);
    signal P_HR_NS241 : unsigned(11 downto 0);
    signal P_HR_NS242 : unsigned(11 downto 0);
    signal P_HR_NS243 : unsigned(11 downto 0);
    signal P_HR_NS244 : unsigned(11 downto 0);
    signal P_HR_NS245 : unsigned(11 downto 0);
    signal P_HR_NS246 : unsigned(11 downto 0);
    signal P_HR_NS247 : unsigned(11 downto 0);
    signal P_HR_NS248 : unsigned(11 downto 0);
    signal P_HR_NS249 : unsigned(11 downto 0);
    signal P_HR_NS250 : unsigned(11 downto 0);
    signal P_HR_NS251 : unsigned(11 downto 0);
    signal P_HR_NS252 : unsigned(11 downto 0);
    signal P_HR_NS253 : unsigned(11 downto 0);
    signal P_HR_NS254 : unsigned(11 downto 0);
    signal P_HR_NS255 : unsigned(11 downto 0);
    signal P_HR_NS256 : unsigned(11 downto 0);
    signal P_HR_NS257 : unsigned(11 downto 0);
    signal P_HR_NS258 : unsigned(11 downto 0);
    signal P_HR_NS259 : unsigned(11 downto 0);
    signal P_HR_NS260 : unsigned(11 downto 0);
    signal P_HR_NS261 : unsigned(11 downto 0);
    signal P_HR_NS262 : unsigned(11 downto 0);
    signal P_HR_NS263 : unsigned(11 downto 0);
    signal P_HR_NS264 : unsigned(11 downto 0);
    signal P_HR_NS265 : unsigned(11 downto 0);
    signal P_HR_NS266 : unsigned(11 downto 0);
    signal P_HR_NS267 : unsigned(11 downto 0);
    signal P_HR_NS268 : unsigned(11 downto 0);
    signal P_HR_NS269 : unsigned(11 downto 0);
    signal P_HR_NS270 : unsigned(11 downto 0);
    signal P_HR_NS271 : unsigned(11 downto 0);
    signal P_HR_NS272 : unsigned(11 downto 0);
    signal P_HR_NS273 : unsigned(11 downto 0);
    signal P_HR_NS274 : unsigned(11 downto 0);
    signal P_HR_NS275 : unsigned(11 downto 0);
    signal P_HR_NS276 : unsigned(11 downto 0);
    signal P_HR_NS277 : unsigned(11 downto 0);
    signal P_HR_NS278 : unsigned(11 downto 0);
    signal P_HR_NS279 : unsigned(11 downto 0);
    signal P_HR_NS280 : unsigned(11 downto 0);
    signal P_HR_NS281 : unsigned(11 downto 0);
    signal P_HR_NS282 : unsigned(11 downto 0);
    signal P_HR_NS283 : unsigned(11 downto 0);
    signal P_HR_NS284 : unsigned(11 downto 0);
    signal P_HR_NS285 : unsigned(11 downto 0);
    signal P_HR_NS286 : unsigned(11 downto 0);
    signal P_HR_NS287 : unsigned(11 downto 0);
    signal P_HR_NS288 : unsigned(11 downto 0);
    signal P_HR_NS289 : unsigned(11 downto 0);
    signal P_HR_NS290 : unsigned(11 downto 0);
    signal P_HR_NS291 : unsigned(11 downto 0);
    signal P_HR_NS292 : unsigned(11 downto 0);
    signal P_HR_NS293 : unsigned(11 downto 0);
    signal P_HR_NS294 : unsigned(11 downto 0);
    signal P_HR_NS295 : unsigned(11 downto 0);
    signal P_HR_NS296 : unsigned(11 downto 0);
    signal P_HR_NS297 : unsigned(11 downto 0);
    signal P_HR_NS298 : unsigned(11 downto 0);
    signal P_HR_NS299 : unsigned(11 downto 0);
    signal P_HR_NS300 : unsigned(11 downto 0);
    signal P_HR_NS301 : unsigned(11 downto 0);
    signal P_HR_NS302 : unsigned(11 downto 0);
    signal P_HR_NS303 : unsigned(11 downto 0);
    signal P_HR_NS304 : unsigned(11 downto 0);
    signal P_HR_NS305 : unsigned(11 downto 0);
    signal P_HR_NS306 : unsigned(11 downto 0);
    signal P_HR_NS307 : unsigned(11 downto 0);
    signal P_HR_NS308 : unsigned(11 downto 0);
    signal P_HR_NS309 : unsigned(11 downto 0);
    signal P_HR_NS310 : unsigned(11 downto 0);
    signal P_HR_NS311 : unsigned(11 downto 0);
    signal P_HR_NS312 : unsigned(11 downto 0);
    signal P_HR_NS313 : unsigned(11 downto 0);
    signal P_HR_NS314 : unsigned(11 downto 0);
    signal P_HR_NS315 : unsigned(11 downto 0);
    signal P_HR_NS316 : unsigned(11 downto 0);
    signal P_HR_NS317 : unsigned(11 downto 0);
    signal P_HR_NS318 : unsigned(11 downto 0);
    signal P_HR_NS319 : unsigned(11 downto 0);
    signal P_HR_NS320 : unsigned(11 downto 0);
    signal P_HR_NS321 : unsigned(11 downto 0);
    signal P_HR_NS322 : unsigned(11 downto 0);
    signal P_HR_NS323 : unsigned(11 downto 0);
    signal P_HR_NS324 : unsigned(11 downto 0);
    signal P_HR_NS325 : unsigned(11 downto 0);
    signal P_HR_NS326 : unsigned(11 downto 0);
    signal P_HR_NS327 : unsigned(11 downto 0);
    signal P_HR_NS328 : unsigned(11 downto 0);
    signal P_HR_NS329 : unsigned(11 downto 0);
    signal P_HR_NS330 : unsigned(11 downto 0);
    signal P_HR_NS331 : unsigned(11 downto 0);
    signal P_HR_NS332 : unsigned(11 downto 0);
    signal P_HR_NS333 : unsigned(11 downto 0);
    signal P_HR_NS334 : unsigned(11 downto 0);
    signal P_HR_NS335 : unsigned(11 downto 0);
    signal P_HR_NS336 : unsigned(11 downto 0);
    signal P_HR_NS337 : unsigned(11 downto 0);
    signal P_HR_NS338 : unsigned(11 downto 0);
    signal P_HR_NS339 : unsigned(11 downto 0);
    signal P_HR_NS340 : unsigned(11 downto 0);
    signal P_HR_NS341 : unsigned(11 downto 0);
    signal P_HR_NS342 : unsigned(11 downto 0);
    signal P_HR_NS343 : unsigned(11 downto 0);
    signal P_HR_NS344 : unsigned(11 downto 0);
    signal P_HR_NS345 : unsigned(11 downto 0);
    signal P_HR_NS346 : unsigned(11 downto 0);
    signal P_HR_NS347 : unsigned(11 downto 0);
    signal P_HR_NS348 : unsigned(11 downto 0);
    signal P_HR_NS349 : unsigned(11 downto 0);
    signal P_HR_NS350 : unsigned(11 downto 0);
    signal P_HR_NS351 : unsigned(11 downto 0);
    signal P_HR_NS352 : unsigned(11 downto 0);
    signal P_HR_NS353 : unsigned(11 downto 0);
    signal P_HR_NS354 : unsigned(11 downto 0);
    signal P_HR_NS355 : unsigned(11 downto 0);
    signal P_HR_NS356 : unsigned(11 downto 0);
    signal P_HR_NS357 : unsigned(11 downto 0);
    signal P_HR_NS358 : unsigned(11 downto 0);
    signal P_HR_NS359 : unsigned(11 downto 0);
    signal P_HR_NS360 : unsigned(11 downto 0);
    signal P_HR_NS361 : unsigned(11 downto 0);
    signal P_HR_NS362 : unsigned(11 downto 0);
    signal P_HR_NS363 : unsigned(11 downto 0);
    signal P_HR_NS364 : unsigned(11 downto 0);
    signal P_HR_NS365 : unsigned(11 downto 0);
    signal P_HR_NS366 : unsigned(11 downto 0);
    signal P_HR_NS367 : unsigned(11 downto 0);
    signal P_HR_NS368 : unsigned(11 downto 0);
    signal P_HR_NS369 : unsigned(11 downto 0);
    signal P_HR_NS370 : unsigned(11 downto 0);
    signal P_HR_NS371 : unsigned(11 downto 0);
    signal P_HR_NS372 : unsigned(11 downto 0);
    signal P_HR_NS373 : unsigned(11 downto 0);
    signal P_HR_NS374 : unsigned(11 downto 0);
    signal P_HR_NS375 : unsigned(11 downto 0);
    signal P_HR_NS376 : unsigned(11 downto 0);
    signal P_HR_NS377 : unsigned(11 downto 0);
    signal P_HR_NS378 : unsigned(11 downto 0);
    signal P_HR_NS379 : unsigned(11 downto 0);
    signal P_HR_NS380 : unsigned(11 downto 0);
    signal P_HR_NS381 : unsigned(11 downto 0);
    signal P_HR_NS382 : unsigned(11 downto 0);
    signal P_HR_NS383 : unsigned(11 downto 0);
    signal P_HR_NS384 : unsigned(11 downto 0);
    signal P_HR_NS385 : unsigned(11 downto 0);
    signal P_HR_NS386 : unsigned(11 downto 0);
    signal P_HR_NS387 : unsigned(11 downto 0);
    signal P_HR_NS388 : unsigned(11 downto 0);
    signal P_HR_NS389 : unsigned(11 downto 0);
    signal P_HR_NS390 : unsigned(11 downto 0);
    signal P_HR_NS391 : unsigned(11 downto 0);
    signal P_HR_NS392 : unsigned(11 downto 0);
    signal P_HR_NS393 : unsigned(11 downto 0);
    signal P_HR_NS394 : unsigned(11 downto 0);
    signal P_HR_NS395 : unsigned(11 downto 0);
    signal P_HR_NS396 : unsigned(11 downto 0);
    signal P_HR_NS397 : unsigned(11 downto 0);
    signal P_HR_NS398 : unsigned(11 downto 0);
    signal P_HR_NS399 : unsigned(11 downto 0);
    signal P_HR_NS400 : unsigned(11 downto 0);
    signal P_HR_NS401 : unsigned(11 downto 0);
    signal P_HR_NS402 : unsigned(11 downto 0);
    signal P_HR_NS403 : unsigned(11 downto 0);
    signal P_HR_NS404 : unsigned(11 downto 0);
    signal P_HR_NS405 : unsigned(11 downto 0);
    signal P_HR_NS406 : unsigned(11 downto 0);
    signal P_HR_NS407 : unsigned(11 downto 0);
    signal P_HR_NS408 : unsigned(11 downto 0);
    signal P_HR_NS409 : unsigned(11 downto 0);
    signal P_HR_NS410 : unsigned(11 downto 0);
    signal P_HR_NS411 : unsigned(11 downto 0);
    signal P_HR_NS412 : unsigned(11 downto 0);
    signal P_HR_NS413 : unsigned(11 downto 0);
    signal P_HR_NS414 : unsigned(11 downto 0);
    signal P_HR_NS415 : unsigned(11 downto 0);
    signal P_HR_NS416 : unsigned(11 downto 0);
    signal P_HR_NS417 : unsigned(11 downto 0);
    signal P_HR_NS418 : unsigned(11 downto 0);
    signal P_HR_NS419 : unsigned(11 downto 0);
    signal P_HR_NS420 : unsigned(11 downto 0);
    signal P_HR_NS421 : unsigned(11 downto 0);
    signal P_HR_NS422 : unsigned(11 downto 0);
    signal P_HR_NS423 : unsigned(11 downto 0);
    signal P_HR_NS424 : unsigned(11 downto 0);
    signal P_HR_NS425 : unsigned(11 downto 0);
    signal P_HR_NS426 : unsigned(11 downto 0);
    signal P_HR_NS427 : unsigned(11 downto 0);
    signal P_HR_NS428 : unsigned(11 downto 0);
    signal P_HR_NS429 : unsigned(11 downto 0);
    signal P_HR_NS430 : unsigned(11 downto 0);
    signal P_HR_NS431 : unsigned(11 downto 0);
    signal P_HR_NS432 : unsigned(11 downto 0);
    signal P_HR_NS433 : unsigned(11 downto 0);
    signal P_HR_NS434 : unsigned(11 downto 0);
    signal P_HR_NS435 : unsigned(11 downto 0);
    signal P_HR_NS436 : unsigned(11 downto 0);
    signal P_HR_NS437 : unsigned(11 downto 0);
    signal P_HR_NS438 : unsigned(11 downto 0);
    signal P_HR_NS439 : unsigned(11 downto 0);
    signal P_HR_NS440 : unsigned(11 downto 0);
    signal P_HR_NS441 : unsigned(11 downto 0);
    signal P_HR_NS442 : unsigned(11 downto 0);
    signal P_HR_NS443 : unsigned(11 downto 0);
    signal P_HR_NS444 : unsigned(11 downto 0);
    signal P_HR_NS445 : unsigned(11 downto 0);
    signal P_HR_NS446 : unsigned(11 downto 0);
    signal P_HR_NS447 : unsigned(11 downto 0);
    signal P_HR_NS448 : unsigned(11 downto 0);
    signal P_HR_NS449 : unsigned(11 downto 0);
    signal P_HR_NS450 : unsigned(11 downto 0);
    signal P_HR_NS451 : unsigned(11 downto 0);
    signal P_HR_NS452 : unsigned(11 downto 0);
    signal P_HR_NS453 : unsigned(11 downto 0);
    signal P_HR_NS454 : unsigned(11 downto 0);
    signal P_HR_NS455 : unsigned(11 downto 0);
    signal P_HR_NS456 : unsigned(11 downto 0);
    signal P_HR_NS457 : unsigned(11 downto 0);
    signal P_HR_NS458 : unsigned(11 downto 0);
    signal P_HR_NS459 : unsigned(11 downto 0);
    signal P_HR_NS460 : unsigned(11 downto 0);
    signal P_HR_NS461 : unsigned(11 downto 0);
    signal P_HR_NS462 : unsigned(11 downto 0);
    signal P_HR_NS463 : unsigned(11 downto 0);
    signal P_HR_NS464 : unsigned(11 downto 0);
    signal P_HR_NS465 : unsigned(11 downto 0);
    signal P_HR_NS466 : unsigned(11 downto 0);
    signal P_HR_NS467 : unsigned(11 downto 0);
    signal P_HR_NS468 : unsigned(11 downto 0);
    signal P_HR_NS469 : unsigned(11 downto 0);
    signal P_HR_NS470 : unsigned(11 downto 0);
    signal P_HR_NS471 : unsigned(11 downto 0);
    signal P_HR_NS472 : unsigned(11 downto 0);
    signal P_HR_NS473 : unsigned(11 downto 0);
    signal P_HR_NS474 : unsigned(11 downto 0);
    signal P_HR_NS475 : unsigned(11 downto 0);
    signal P_HR_NS476 : unsigned(11 downto 0);
    signal P_HR_NS477 : unsigned(11 downto 0);
    signal P_HR_NS478 : unsigned(11 downto 0);
    signal P_HR_NS479 : unsigned(11 downto 0);
    signal P_HR_NS480 : unsigned(11 downto 0);
    signal P_HR_NS481 : unsigned(11 downto 0);
    signal P_HR_NS482 : unsigned(11 downto 0);
    signal P_HR_NS483 : unsigned(11 downto 0);
    signal P_HR_NS484 : unsigned(11 downto 0);
    signal P_HR_NS485 : unsigned(11 downto 0);
    signal P_HR_NS486 : unsigned(11 downto 0);
    signal P_HR_NS487 : unsigned(11 downto 0);
    signal P_HR_NS488 : unsigned(11 downto 0);
    signal P_HR_NS489 : unsigned(11 downto 0);
    signal P_HR_NS490 : unsigned(11 downto 0);
    signal P_HR_NS491 : unsigned(11 downto 0);
    signal P_HR_NS492 : unsigned(11 downto 0);
    signal P_HR_NS493 : unsigned(11 downto 0);
    signal P_HR_NS494 : unsigned(11 downto 0);
    signal P_HR_NS495 : unsigned(11 downto 0);
    signal P_HR_NS496 : unsigned(11 downto 0);
    signal P_HR_NS497 : unsigned(11 downto 0);
    signal P_HR_NS498 : unsigned(11 downto 0);
    signal P_HR_NS499 : unsigned(11 downto 0);
    signal P_HR_NS500 : unsigned(11 downto 0);
    signal P_HR_NS501 : unsigned(11 downto 0);
    signal P_HR_NS502 : unsigned(11 downto 0);
    signal P_HR_NS503 : unsigned(11 downto 0);
    signal P_HR_NS504 : unsigned(11 downto 0);
    signal P_HR_NS505 : unsigned(11 downto 0);
    signal P_HR_NS506 : unsigned(11 downto 0);
    signal P_HR_NS507 : unsigned(11 downto 0);
    signal P_HR_NS508 : unsigned(11 downto 0);
    signal P_HR_NS509 : unsigned(11 downto 0);
    signal P_HR_NS510 : unsigned(11 downto 0);
    signal P_HR_NS511 : unsigned(11 downto 0);
    signal P_HR_NS512 : unsigned(11 downto 0);
    signal P_HR_NS513 : unsigned(11 downto 0);
    signal P_HR_NS514 : unsigned(11 downto 0);
    signal P_HR_NS515 : unsigned(11 downto 0);
    signal P_HR_NS516 : unsigned(11 downto 0);
    signal P_HR_NS517 : unsigned(11 downto 0);
    signal P_HR_NS518 : unsigned(11 downto 0);
    signal P_HR_NS519 : unsigned(11 downto 0);
    signal P_HR_NS520 : unsigned(11 downto 0);
    signal P_HR_NS521 : unsigned(11 downto 0);
    signal P_HR_NS522 : unsigned(11 downto 0);
    signal P_HR_NS523 : unsigned(11 downto 0);
    signal P_HR_NS524 : unsigned(11 downto 0);
    signal P_HR_NS525 : unsigned(11 downto 0);
    signal P_HR_NS526 : unsigned(11 downto 0);
    signal P_HR_NS527 : unsigned(11 downto 0);
    signal P_HR_NS528 : unsigned(11 downto 0);
    signal P_HR_NS529 : unsigned(11 downto 0);
    signal P_HR_NS530 : unsigned(11 downto 0);
    signal P_HR_NS531 : unsigned(11 downto 0);
    signal P_HR_NS532 : unsigned(11 downto 0);
    signal P_HR_NS533 : unsigned(11 downto 0);
    signal P_HR_NS534 : unsigned(11 downto 0);
    signal P_HR_NS535 : unsigned(11 downto 0);
    signal P_HR_NS536 : unsigned(11 downto 0);
    signal P_HR_NS537 : unsigned(11 downto 0);
    signal P_HR_NS538 : unsigned(11 downto 0);
    signal P_HR_NS539 : unsigned(11 downto 0);
    signal P_HR_NS540 : unsigned(11 downto 0);
    signal P_HR_NS541 : unsigned(11 downto 0);
    signal P_HR_NS542 : unsigned(11 downto 0);
    signal P_HR_NS543 : unsigned(11 downto 0);
    signal P_HR_NS544 : unsigned(11 downto 0);
    signal P_HR_NS545 : unsigned(11 downto 0);
    signal P_HR_NS546 : unsigned(11 downto 0);
    signal P_HR_NS547 : unsigned(11 downto 0);
    signal P_HR_NS548 : unsigned(11 downto 0);
    signal P_HR_NS549 : unsigned(11 downto 0);
    signal P_HR_NS550 : unsigned(11 downto 0);
    signal P_HR_NS551 : unsigned(11 downto 0);
    signal P_HR_NS552 : unsigned(11 downto 0);
    signal P_HR_NS553 : unsigned(11 downto 0);
    signal P_HR_NS554 : unsigned(11 downto 0);
    signal P_HR_NS555 : unsigned(11 downto 0);
    signal P_HR_NS556 : unsigned(11 downto 0);
    signal P_HR_NS557 : unsigned(11 downto 0);
    signal P_HR_NS558 : unsigned(11 downto 0);
    signal P_HR_NS559 : unsigned(11 downto 0);
    signal P_HR_NS560 : unsigned(11 downto 0);
    signal P_HR_NS561 : unsigned(11 downto 0);
    signal P_HR_NS562 : unsigned(11 downto 0);
    signal P_HR_NS563 : unsigned(11 downto 0);
    signal P_HR_NS564 : unsigned(11 downto 0);
    signal P_HR_NS565 : unsigned(11 downto 0);
    signal P_HR_NS566 : unsigned(11 downto 0);
    signal P_HR_NS567 : unsigned(11 downto 0);
    signal P_HR_NS568 : unsigned(11 downto 0);
    signal P_HR_NS569 : unsigned(11 downto 0);
    signal P_HR_NS570 : unsigned(11 downto 0);
    signal P_HR_NS571 : unsigned(11 downto 0);
    signal P_HR_NS572 : unsigned(11 downto 0);
    signal P_HR_NS573 : unsigned(11 downto 0);
    signal P_HR_NS574 : unsigned(11 downto 0);
    signal P_HR_NS575 : unsigned(11 downto 0);
    signal P_HR_NS576 : unsigned(11 downto 0);
    signal P_HR_NS577 : unsigned(11 downto 0);
    signal P_HR_NS578 : unsigned(11 downto 0);
    signal P_HR_NS579 : unsigned(11 downto 0);
    signal P_HR_NS580 : unsigned(11 downto 0);
    signal P_HR_NS581 : unsigned(11 downto 0);
    signal P_HR_NS582 : unsigned(11 downto 0);
    signal P_HR_NS583 : unsigned(11 downto 0);
    signal P_HR_NS584 : unsigned(11 downto 0);
    signal P_HR_NS585 : unsigned(11 downto 0);
    signal P_HR_NS586 : unsigned(11 downto 0);
    signal P_HR_NS587 : unsigned(11 downto 0);
    signal P_HR_NS588 : unsigned(11 downto 0);
    signal P_HR_NS589 : unsigned(11 downto 0);
    signal P_HR_NS590 : unsigned(11 downto 0);
    signal P_HR_NS591 : unsigned(11 downto 0);
    signal P_HR_NS592 : unsigned(11 downto 0);
    signal P_HR_NS593 : unsigned(11 downto 0);
    signal P_HR_NS594 : unsigned(11 downto 0);
    signal P_HR_NS595 : unsigned(11 downto 0);
    signal P_HR_NS596 : unsigned(11 downto 0);
    signal P_HR_NS597 : unsigned(11 downto 0);
    signal P_HR_NS598 : unsigned(11 downto 0);
    signal P_HR_NS599 : unsigned(11 downto 0);
    signal P_HR_NS600 : unsigned(11 downto 0);
    signal P_HR_NS601 : unsigned(11 downto 0);
    signal P_HR_NS602 : unsigned(11 downto 0);
    signal P_HR_NS603 : unsigned(11 downto 0);
    signal P_HR_NS604 : unsigned(11 downto 0);
    signal P_HR_NS605 : unsigned(11 downto 0);
    signal P_HR_NS606 : unsigned(11 downto 0);
    signal P_HR_NS607 : unsigned(11 downto 0);
    signal P_HR_NS608 : unsigned(11 downto 0);
    signal P_HR_NS609 : unsigned(11 downto 0);
    signal P_HR_NS610 : unsigned(11 downto 0);
    signal P_HR_NS611 : unsigned(11 downto 0);
    signal P_HR_NS612 : unsigned(11 downto 0);
    signal P_HR_NS613 : unsigned(11 downto 0);
    signal P_HR_NS614 : unsigned(11 downto 0);
    signal P_HR_NS615 : unsigned(11 downto 0);
    signal P_HR_NS616 : unsigned(11 downto 0);
    signal P_HR_NS617 : unsigned(11 downto 0);
    signal P_HR_NS618 : unsigned(11 downto 0);
    signal P_HR_NS619 : unsigned(11 downto 0);
    signal P_HR_NS620 : unsigned(11 downto 0);
    signal P_HR_NS621 : unsigned(11 downto 0);
    signal P_HR_NS622 : unsigned(11 downto 0);
    signal P_HR_NS623 : unsigned(11 downto 0);
    signal P_HR_NS624 : unsigned(11 downto 0);
    signal P_HR_NS625 : unsigned(11 downto 0);
    signal P_HR_NS626 : unsigned(11 downto 0);
    signal P_HR_NS627 : unsigned(11 downto 0);
    signal P_HR_NS628 : unsigned(11 downto 0);
    signal P_HR_NS629 : unsigned(11 downto 0);
    signal P_HR_NS630 : unsigned(11 downto 0);
    signal P_HR_NS631 : unsigned(11 downto 0);
    signal P_HR_NS632 : unsigned(11 downto 0);
    signal P_HR_NS633 : unsigned(11 downto 0);
    signal P_HR_NS634 : unsigned(11 downto 0);
    signal P_HR_NS635 : unsigned(11 downto 0);
    signal P_HR_NS636 : unsigned(11 downto 0);
    signal P_HR_NS637 : unsigned(11 downto 0);
    signal P_HR_NS638 : unsigned(11 downto 0);
    signal P_HR_NS639 : unsigned(11 downto 0);
    signal P_HR_NS640 : unsigned(11 downto 0);
    signal P_HR_NS641 : unsigned(11 downto 0);
    signal P_HR_NS642 : unsigned(11 downto 0);
    signal P_HR_NS643 : unsigned(11 downto 0);
    signal P_HR_NS644 : unsigned(11 downto 0);
    signal P_HR_NS645 : unsigned(11 downto 0);
    signal P_HR_NS646 : unsigned(11 downto 0);
    signal P_HR_NS647 : unsigned(11 downto 0);
    signal P_HR_NS648 : unsigned(11 downto 0);
    signal P_HR_NS649 : unsigned(11 downto 0);
    signal P_HR_NS650 : unsigned(11 downto 0);
    signal P_HR_NS651 : unsigned(11 downto 0);
    signal P_HR_NS652 : unsigned(11 downto 0);
    signal P_HR_NS653 : unsigned(11 downto 0);
    signal P_HR_NS654 : unsigned(11 downto 0);
    signal P_HR_NS655 : unsigned(11 downto 0);
    signal P_HR_NS656 : unsigned(11 downto 0);
    signal P_HR_NS657 : unsigned(11 downto 0);
    signal P_HR_NS658 : unsigned(11 downto 0);
    signal P_HR_NS659 : unsigned(11 downto 0);
    signal P_HR_NS660 : unsigned(11 downto 0);
    signal P_HR_NS661 : unsigned(11 downto 0);
    signal P_HR_NS662 : unsigned(11 downto 0);
    signal P_HR_NS663 : unsigned(11 downto 0);
    signal P_HR_NS664 : unsigned(11 downto 0);
    signal P_HR_NS665 : unsigned(11 downto 0);
    signal P_HR_NS666 : unsigned(11 downto 0);
    signal P_HR_NS667 : unsigned(11 downto 0);
    signal P_HR_NS668 : unsigned(11 downto 0);
    signal P_HR_NS669 : unsigned(11 downto 0);
    signal P_HR_NS670 : unsigned(11 downto 0);
    signal P_HR_NS671 : unsigned(11 downto 0);
    signal P_HR_NS672 : unsigned(11 downto 0);
    signal P_HR_NS673 : unsigned(11 downto 0);
    signal P_HR_NS674 : unsigned(11 downto 0);
    signal P_HR_NS675 : unsigned(11 downto 0);
    signal P_HR_NS676 : unsigned(11 downto 0);
    signal P_HR_NS677 : unsigned(11 downto 0);
    signal P_HR_NS678 : unsigned(11 downto 0);
    signal P_HR_NS679 : unsigned(11 downto 0);
    signal P_HR_NS680 : unsigned(11 downto 0);
    signal P_HR_NS681 : unsigned(11 downto 0);
    signal P_HR_NS682 : unsigned(11 downto 0);
    signal P_HR_NS683 : unsigned(11 downto 0);
    signal P_HR_NS684 : unsigned(11 downto 0);
    signal P_HR_NS685 : unsigned(11 downto 0);
    signal P_HR_NS686 : unsigned(11 downto 0);
    signal P_HR_NS687 : unsigned(11 downto 0);
    signal P_HR_NS688 : unsigned(11 downto 0);
    signal P_HR_NS689 : unsigned(11 downto 0);
    signal P_HR_NS690 : unsigned(11 downto 0);
    signal P_HR_NS691 : unsigned(11 downto 0);
    signal P_HR_NS692 : unsigned(11 downto 0);
    signal P_HR_NS693 : unsigned(11 downto 0);
    signal P_HR_NS694 : unsigned(11 downto 0);
    signal P_HR_NS695 : unsigned(11 downto 0);
    signal P_HR_NS696 : unsigned(11 downto 0);
    signal P_HR_NS697 : unsigned(11 downto 0);
    signal P_HR_NS698 : unsigned(11 downto 0);
    signal P_HR_NS699 : unsigned(11 downto 0);
    signal P_HR_NS700 : unsigned(11 downto 0);
    signal P_HR_NS701 : unsigned(11 downto 0);
    signal P_HR_NS702 : unsigned(11 downto 0);
    signal P_HR_NS703 : unsigned(11 downto 0);
    signal P_HR_NS704 : unsigned(11 downto 0);
    signal P_HR_NS705 : unsigned(11 downto 0);
    signal P_HR_NS706 : unsigned(11 downto 0);
    signal P_HR_NS707 : unsigned(11 downto 0);
    signal P_HR_NS708 : unsigned(11 downto 0);
    signal P_HR_NS709 : unsigned(11 downto 0);
    signal P_HR_NS710 : unsigned(11 downto 0);
    signal P_HR_NS711 : unsigned(11 downto 0);
    signal P_HR_NS712 : unsigned(11 downto 0);
    signal P_HR_NS713 : unsigned(11 downto 0);
    signal P_HR_NS714 : unsigned(11 downto 0);
    signal P_HR_NS715 : unsigned(11 downto 0);
    signal P_HR_NS716 : unsigned(11 downto 0);
    signal P_HR_NS717 : unsigned(11 downto 0);
    signal P_HR_NS718 : unsigned(11 downto 0);
    signal P_HR_NS719 : unsigned(11 downto 0);
    signal P_HR_NS720 : unsigned(11 downto 0);
    signal P_HR_NS721 : unsigned(11 downto 0);
    signal P_HR_NS722 : unsigned(11 downto 0);
    signal P_HR_NS723 : unsigned(11 downto 0);
    signal P_HR_NS724 : unsigned(11 downto 0);
    signal P_HR_NS725 : unsigned(11 downto 0);
    signal P_HR_NS726 : unsigned(11 downto 0);
		
    signal P_EDA_NS1 : unsigned(11 downto 0);
    signal P_EDA_NS2 : unsigned(11 downto 0);
    signal P_EDA_NS3 : unsigned(11 downto 0);
    signal P_EDA_NS4 : unsigned(11 downto 0);
    signal P_EDA_NS5 : unsigned(11 downto 0);
    signal P_EDA_NS6 : unsigned(11 downto 0);
    signal P_EDA_NS7 : unsigned(11 downto 0);
    signal P_EDA_NS8 : unsigned(11 downto 0);
    signal P_EDA_NS9 : unsigned(11 downto 0);
    signal P_EDA_NS10 : unsigned(11 downto 0);
    signal P_EDA_NS11 : unsigned(11 downto 0);
    signal P_EDA_NS12 : unsigned(11 downto 0);
    signal P_EDA_NS13 : unsigned(11 downto 0);
    signal P_EDA_NS14 : unsigned(11 downto 0);
    signal P_EDA_NS15 : unsigned(11 downto 0);
    signal P_EDA_NS16 : unsigned(11 downto 0);
    signal P_EDA_NS17 : unsigned(11 downto 0);
    signal P_EDA_NS18 : unsigned(11 downto 0);
    signal P_EDA_NS19 : unsigned(11 downto 0);
    signal P_EDA_NS20 : unsigned(11 downto 0);
    signal P_EDA_NS21 : unsigned(11 downto 0);
    signal P_EDA_NS22 : unsigned(11 downto 0);
    signal P_EDA_NS23 : unsigned(11 downto 0);
    signal P_EDA_NS24 : unsigned(11 downto 0);
    signal P_EDA_NS25 : unsigned(11 downto 0);
    signal P_EDA_NS26 : unsigned(11 downto 0);
    signal P_EDA_NS27 : unsigned(11 downto 0);
    signal P_EDA_NS28 : unsigned(11 downto 0);
    signal P_EDA_NS29 : unsigned(11 downto 0);
    signal P_EDA_NS30 : unsigned(11 downto 0);
    signal P_EDA_NS31 : unsigned(11 downto 0);
    signal P_EDA_NS32 : unsigned(11 downto 0);
    signal P_EDA_NS33 : unsigned(11 downto 0);
    signal P_EDA_NS34 : unsigned(11 downto 0);
    signal P_EDA_NS35 : unsigned(11 downto 0);
    signal P_EDA_NS36 : unsigned(11 downto 0);
    signal P_EDA_NS37 : unsigned(11 downto 0);
    signal P_EDA_NS38 : unsigned(11 downto 0);
    signal P_EDA_NS39 : unsigned(11 downto 0);
    signal P_EDA_NS40 : unsigned(11 downto 0);
    signal P_EDA_NS41 : unsigned(11 downto 0);
    signal P_EDA_NS42 : unsigned(11 downto 0);
    signal P_EDA_NS43 : unsigned(11 downto 0);
    signal P_EDA_NS44 : unsigned(11 downto 0);
    signal P_EDA_NS45 : unsigned(11 downto 0);
    signal P_EDA_NS46 : unsigned(11 downto 0);
    signal P_EDA_NS47 : unsigned(11 downto 0);
    signal P_EDA_NS48 : unsigned(11 downto 0);
    signal P_EDA_NS49 : unsigned(11 downto 0);
    signal P_EDA_NS50 : unsigned(11 downto 0);
    signal P_EDA_NS51 : unsigned(11 downto 0);
    signal P_EDA_NS52 : unsigned(11 downto 0);
    signal P_EDA_NS53 : unsigned(11 downto 0);
    signal P_EDA_NS54 : unsigned(11 downto 0);
    signal P_EDA_NS55 : unsigned(11 downto 0);
    signal P_EDA_NS56 : unsigned(11 downto 0);
    signal P_EDA_NS57 : unsigned(11 downto 0);
    signal P_EDA_NS58 : unsigned(11 downto 0);
    signal P_EDA_NS59 : unsigned(11 downto 0);
    signal P_EDA_NS60 : unsigned(11 downto 0);
    signal P_EDA_NS61 : unsigned(11 downto 0);
    signal P_EDA_NS62 : unsigned(11 downto 0);
    signal P_EDA_NS63 : unsigned(11 downto 0);
    signal P_EDA_NS64 : unsigned(11 downto 0);
    signal P_EDA_NS65 : unsigned(11 downto 0);
    signal P_EDA_NS66 : unsigned(11 downto 0);
    signal P_EDA_NS67 : unsigned(11 downto 0);
    signal P_EDA_NS68 : unsigned(11 downto 0);
    signal P_EDA_NS69 : unsigned(11 downto 0);
    signal P_EDA_NS70 : unsigned(11 downto 0);
    signal P_EDA_NS71 : unsigned(11 downto 0);
    signal P_EDA_NS72 : unsigned(11 downto 0);
    signal P_EDA_NS73 : unsigned(11 downto 0);
    signal P_EDA_NS74 : unsigned(11 downto 0);
    signal P_EDA_NS75 : unsigned(11 downto 0);
    signal P_EDA_NS76 : unsigned(11 downto 0);
    signal P_EDA_NS77 : unsigned(11 downto 0);
    signal P_EDA_NS78 : unsigned(11 downto 0);
    signal P_EDA_NS79 : unsigned(11 downto 0);
    signal P_EDA_NS80 : unsigned(11 downto 0);
    signal P_EDA_NS81 : unsigned(11 downto 0);
    signal P_EDA_NS82 : unsigned(11 downto 0);
    signal P_EDA_NS83 : unsigned(11 downto 0);
    signal P_EDA_NS84 : unsigned(11 downto 0);
    signal P_EDA_NS85 : unsigned(11 downto 0);
    signal P_EDA_NS86 : unsigned(11 downto 0);
    signal P_EDA_NS87 : unsigned(11 downto 0);
    signal P_EDA_NS88 : unsigned(11 downto 0);
    signal P_EDA_NS89 : unsigned(11 downto 0);
    signal P_EDA_NS90 : unsigned(11 downto 0);
    signal P_EDA_NS91 : unsigned(11 downto 0);
    signal P_EDA_NS92 : unsigned(11 downto 0);
    signal P_EDA_NS93 : unsigned(11 downto 0);
    signal P_EDA_NS94 : unsigned(11 downto 0);
    signal P_EDA_NS95 : unsigned(11 downto 0);
    signal P_EDA_NS96 : unsigned(11 downto 0);
    signal P_EDA_NS97 : unsigned(11 downto 0);
    signal P_EDA_NS98 : unsigned(11 downto 0);
    signal P_EDA_NS99 : unsigned(11 downto 0);
    signal P_EDA_NS100 : unsigned(11 downto 0);
    signal P_EDA_NS101 : unsigned(11 downto 0);
    signal P_EDA_NS102 : unsigned(11 downto 0);
    signal P_EDA_NS103 : unsigned(11 downto 0);
    signal P_EDA_NS104 : unsigned(11 downto 0);
    signal P_EDA_NS105 : unsigned(11 downto 0);
    signal P_EDA_NS106 : unsigned(11 downto 0);
    signal P_EDA_NS107 : unsigned(11 downto 0);
    signal P_EDA_NS108 : unsigned(11 downto 0);
    signal P_EDA_NS109 : unsigned(11 downto 0);
    signal P_EDA_NS110 : unsigned(11 downto 0);
	
	signal P_TEMP_S : unsigned(11 downto 0);
	signal P_TEMP_NS : unsigned(11 downto 0);
	
	signal P_EDA_S : unsigned(11 downto 0);
	signal P_EDA_NS : unsigned(11 downto 0);
	
	signal P_HR_S : unsigned(11 downto 0);
	signal P_HR_NS : unsigned(11 downto 0);
	
	signal stress_score : unsigned(47 downto 0);
	signal not_stress_score : unsigned(48 downto 0);
	
	type type_state is (NORMAL, TRAINING_S, TRAINING_NS);
	attribute enum_encoding : string;
	attribute enum_encoding of type_state : type is "00 01 11";
	
	signal state, next_state: type_state;
	
	-- constants
    constant P_STRESS : unsigned(11 downto 0) := "011111010000"; -- 20
	constant P_NOT_STRESS : unsigned(12 downto 0) := "1111101000000"; -- 80
	constant T_STRESS : unsigned(5 downto 0) := "001000";
	constant T_N_STRESS : unsigned(5 downto 0) := "000001";
	
	--constant P_STRESS : unsigned(12 downto 0) := "1001110001000"; 
	--constant P_NOT_STRESS : unsigned(12 downto 0) := "1001110001000";
	
begin
	
	process(clk, rst) --state transition
	begin
		if (rst = '1') then
			state <= NORMAL;
		elsif (rising_edge(clk)) then
			state <= next_state;
		end if;
	end process;
	
	process(state, s1) -- combinational state assignment
	begin
		case state is
			when NORMAL =>
				if s1 = "01" then
					next_state <= TRAINING_S;
				elsif s1 = "11" then
					next_state <= TRAINING_NS;
				else
					next_state <= NORMAL;
				end if;
			when TRAINING_S =>
				if s1 = "01" then
					next_state <= TRAINING_S;
				elsif s1 = "11" then
					next_state <= TRAINING_NS;
				else
					next_state <= NORMAL;
				end if;
			when TRAINING_NS =>
				if s1 = "01" then
					next_state <= TRAINING_S;
				elsif s1 = "11" then
					next_state <= TRAINING_NS;
				else
					next_state <= NORMAL;
				end if;
			when others => null;
		end case;
	end process;
	
	-- should expect status = 11 when in training mode
	process(clk,rst) -- output block
	begin
		if (rst = '1') then
			status <= "00";
		elsif (rising_edge(clk)) then
			if stress_score < not_stress_score then
				status <= "01"; -- not stressed
			elsif stress_score > not_stress_score then
				status <= "10"; -- stressed
			elsif stress_score = not_stress_score then
				status <= "11"; -- rare, equality
			else
				status <= "00";
			end if;

		end if;	
	end process;	
	

	process(clk, rst) -- stress score
	begin
		if (rst = '1') then
		-- reset logic
        P_TEMP_S1 <= (others => '0');
        P_TEMP_S2 <= (others => '0');
        P_TEMP_S3 <= (others => '0');
        P_TEMP_S4 <= (others => '0');
        P_TEMP_S5 <= (others => '0');
        P_TEMP_S6 <= (others => '0');
        P_TEMP_S7 <= (others => '0');
        P_TEMP_S8 <= (others => '0');
        P_TEMP_S9 <= (others => '0');
        P_TEMP_S10 <= (others => '0');
        P_TEMP_S11 <= (others => '0');
        P_TEMP_S12 <= (others => '0');
        P_TEMP_S13 <= (others => '0');
        P_TEMP_S14 <= (others => '0');
        P_TEMP_S15 <= (others => '0');
        P_TEMP_S16 <= (others => '0');
        P_TEMP_S17 <= (others => '0');
        P_TEMP_S18 <= (others => '0');
        P_TEMP_S19 <= (others => '0');
        P_TEMP_S20 <= (others => '0');
        P_TEMP_S21 <= (others => '0');
        P_TEMP_S22 <= (others => '0');
        P_TEMP_S23 <= (others => '0');
        P_TEMP_S24 <= (others => '0');
        P_TEMP_S25 <= (others => '0');
        P_TEMP_S26 <= (others => '0');
        P_TEMP_S27 <= (others => '0');
        P_TEMP_S28 <= (others => '0');
        P_TEMP_S29 <= (others => '0');
        P_TEMP_S30 <= (others => '0');
        P_TEMP_S31 <= (others => '0');
        P_TEMP_S32 <= (others => '0');
        P_TEMP_S33 <= (others => '0');
        P_TEMP_S34 <= (others => '0');
        P_TEMP_S35 <= (others => '0');
        P_TEMP_S36 <= (others => '0');
        P_TEMP_S37 <= (others => '0');
        P_TEMP_S38 <= (others => '0');
        P_TEMP_S39 <= (others => '0');
        P_TEMP_S40 <= (others => '0');
			
        P_EDA_S1 <= (others => '0');
        P_EDA_S2 <= (others => '0');
        P_EDA_S3 <= (others => '0');
        P_EDA_S4 <= (others => '0');
        P_EDA_S5 <= (others => '0');
        P_EDA_S6 <= (others => '0');
        P_EDA_S7 <= (others => '0');
        P_EDA_S8 <= (others => '0');
        P_EDA_S9 <= (others => '0');
        P_EDA_S10 <= (others => '0');
        P_EDA_S11 <= (others => '0');
        P_EDA_S12 <= (others => '0');
        P_EDA_S13 <= (others => '0');
        P_EDA_S14 <= (others => '0');
        P_EDA_S15 <= (others => '0');
        P_EDA_S16 <= (others => '0');
        P_EDA_S17 <= (others => '0');
        P_EDA_S18 <= (others => '0');
        P_EDA_S19 <= (others => '0');
        P_EDA_S20 <= (others => '0');
        P_EDA_S21 <= (others => '0');
        P_EDA_S22 <= (others => '0');
        P_EDA_S23 <= (others => '0');
        P_EDA_S24 <= (others => '0');
        P_EDA_S25 <= (others => '0');
        P_EDA_S26 <= (others => '0');
        P_EDA_S27 <= (others => '0');
        P_EDA_S28 <= (others => '0');
        P_EDA_S29 <= (others => '0');
        P_EDA_S30 <= (others => '0');
        P_EDA_S31 <= (others => '0');
        P_EDA_S32 <= (others => '0');
        P_EDA_S33 <= (others => '0');
        P_EDA_S34 <= (others => '0');
        P_EDA_S35 <= (others => '0');
        P_EDA_S36 <= (others => '0');
        P_EDA_S37 <= (others => '0');
        P_EDA_S38 <= (others => '0');
        P_EDA_S39 <= (others => '0');
        P_EDA_S40 <= (others => '0');
        P_EDA_S41 <= (others => '0');
        P_EDA_S42 <= (others => '0');
        P_EDA_S43 <= (others => '0');
        P_EDA_S44 <= (others => '0');
        P_EDA_S45 <= (others => '0');
        P_EDA_S46 <= (others => '0');
        P_EDA_S47 <= (others => '0');
        P_EDA_S48 <= (others => '0');
        P_EDA_S49 <= (others => '0');
        P_EDA_S50 <= (others => '0');
        P_EDA_S51 <= (others => '0');
        P_EDA_S52 <= (others => '0');
        P_EDA_S53 <= (others => '0');
        P_EDA_S54 <= (others => '0');
        P_EDA_S55 <= (others => '0');
        P_EDA_S56 <= (others => '0');
        P_EDA_S57 <= (others => '0');
        P_EDA_S58 <= (others => '0');
        P_EDA_S59 <= (others => '0');
        P_EDA_S60 <= (others => '0');
        P_EDA_S61 <= (others => '0');
        P_EDA_S62 <= (others => '0');
        P_EDA_S63 <= (others => '0');
        P_EDA_S64 <= (others => '0');
        P_EDA_S65 <= (others => '0');
        P_EDA_S66 <= (others => '0');
        P_EDA_S67 <= (others => '0');
        P_EDA_S68 <= (others => '0');
        P_EDA_S69 <= (others => '0');
        P_EDA_S70 <= (others => '0');
        P_EDA_S71 <= (others => '0');
        P_EDA_S72 <= (others => '0');
        P_EDA_S73 <= (others => '0');
        P_EDA_S74 <= (others => '0');
        P_EDA_S75 <= (others => '0');
        P_EDA_S76 <= (others => '0');
        P_EDA_S77 <= (others => '0');
        P_EDA_S78 <= (others => '0');
        P_EDA_S79 <= (others => '0');
        P_EDA_S80 <= (others => '0');
        P_EDA_S81 <= (others => '0');
        P_EDA_S82 <= (others => '0');
        P_EDA_S83 <= (others => '0');
        P_EDA_S84 <= (others => '0');
        P_EDA_S85 <= (others => '0');
        P_EDA_S86 <= (others => '0');
        P_EDA_S87 <= (others => '0');
        P_EDA_S88 <= (others => '0');
        P_EDA_S89 <= (others => '0');
        P_EDA_S90 <= (others => '0');
        P_EDA_S91 <= (others => '0');
        P_EDA_S92 <= (others => '0');
        P_EDA_S93 <= (others => '0');
        P_EDA_S94 <= (others => '0');
        P_EDA_S95 <= (others => '0');
        P_EDA_S96 <= (others => '0');
        P_EDA_S97 <= (others => '0');
        P_EDA_S98 <= (others => '0');
        P_EDA_S99 <= (others => '0');
        P_EDA_S100 <= (others => '0');
        P_EDA_S101 <= (others => '0');
        P_EDA_S102 <= (others => '0');
        P_EDA_S103 <= (others => '0');
        P_EDA_S104 <= (others => '0');
        P_EDA_S105 <= (others => '0');
        P_EDA_S106 <= (others => '0');
        P_EDA_S107 <= (others => '0');
        P_EDA_S108 <= (others => '0');
        P_EDA_S109 <= (others => '0');
        P_EDA_S110 <= (others => '0');
        P_EDA_S111 <= (others => '0');
        P_EDA_S112 <= (others => '0');
        P_EDA_S113 <= (others => '0');
        P_EDA_S114 <= (others => '0');
        P_EDA_S115 <= (others => '0');
        P_EDA_S116 <= (others => '0');
        P_EDA_S117 <= (others => '0');
        P_EDA_S118 <= (others => '0');
        P_EDA_S119 <= (others => '0');
        P_EDA_S120 <= (others => '0');
        P_EDA_S121 <= (others => '0');
        P_EDA_S122 <= (others => '0');
        P_EDA_S123 <= (others => '0');
        P_EDA_S124 <= (others => '0');
        P_EDA_S125 <= (others => '0');
        P_EDA_S126 <= (others => '0');
        P_EDA_S127 <= (others => '0');
        P_EDA_S128 <= (others => '0');
        P_EDA_S129 <= (others => '0');
        P_EDA_S130 <= (others => '0');
			
        P_HR_S1 <= (others => '0');
        P_HR_S2 <= (others => '0');
        P_HR_S3 <= (others => '0');
        P_HR_S4 <= (others => '0');
        P_HR_S5 <= (others => '0');
        P_HR_S6 <= (others => '0');
        P_HR_S7 <= (others => '0');
        P_HR_S8 <= (others => '0');
        P_HR_S9 <= (others => '0');
        P_HR_S10 <= (others => '0');
        P_HR_S11 <= (others => '0');
        P_HR_S12 <= (others => '0');
        P_HR_S13 <= (others => '0');
        P_HR_S14 <= (others => '0');
        P_HR_S15 <= (others => '0');
        P_HR_S16 <= (others => '0');
        P_HR_S17 <= (others => '0');
        P_HR_S18 <= (others => '0');
        P_HR_S19 <= (others => '0');
        P_HR_S20 <= (others => '0');
        P_HR_S21 <= (others => '0');
        P_HR_S22 <= (others => '0');
        P_HR_S23 <= (others => '0');
        P_HR_S24 <= (others => '0');
        P_HR_S25 <= (others => '0');
        P_HR_S26 <= (others => '0');
        P_HR_S27 <= (others => '0');
        P_HR_S28 <= (others => '0');
        P_HR_S29 <= (others => '0');
        P_HR_S30 <= (others => '0');
        P_HR_S31 <= (others => '0');
        P_HR_S32 <= (others => '0');
        P_HR_S33 <= (others => '0');
        P_HR_S34 <= (others => '0');
        P_HR_S35 <= (others => '0');
        P_HR_S36 <= (others => '0');
        P_HR_S37 <= (others => '0');
        P_HR_S38 <= (others => '0');
        P_HR_S39 <= (others => '0');
        P_HR_S40 <= (others => '0');
        P_HR_S41 <= (others => '0');
        P_HR_S42 <= (others => '0');
        P_HR_S43 <= (others => '0');
        P_HR_S44 <= (others => '0');
        P_HR_S45 <= (others => '0');
        P_HR_S46 <= (others => '0');
        P_HR_S47 <= (others => '0');
        P_HR_S48 <= (others => '0');
        P_HR_S49 <= (others => '0');
        P_HR_S50 <= (others => '0');
        P_HR_S51 <= (others => '0');
        P_HR_S52 <= (others => '0');
        P_HR_S53 <= (others => '0');
        P_HR_S54 <= (others => '0');
        P_HR_S55 <= (others => '0');
        P_HR_S56 <= (others => '0');
        P_HR_S57 <= (others => '0');
        P_HR_S58 <= (others => '0');
        P_HR_S59 <= (others => '0');
        P_HR_S60 <= (others => '0');
        P_HR_S61 <= (others => '0');
        P_HR_S62 <= (others => '0');
        P_HR_S63 <= (others => '0');
        P_HR_S64 <= (others => '0');
        P_HR_S65 <= (others => '0');
        P_HR_S66 <= (others => '0');
        P_HR_S67 <= (others => '0');
        P_HR_S68 <= (others => '0');
        P_HR_S69 <= (others => '0');
        P_HR_S70 <= (others => '0');
        P_HR_S71 <= (others => '0');
        P_HR_S72 <= (others => '0');
        P_HR_S73 <= (others => '0');
        P_HR_S74 <= (others => '0');
        P_HR_S75 <= (others => '0');
        P_HR_S76 <= (others => '0');
        P_HR_S77 <= (others => '0');
        P_HR_S78 <= (others => '0');
        P_HR_S79 <= (others => '0');
        P_HR_S80 <= (others => '0');
        P_HR_S81 <= (others => '0');
        P_HR_S82 <= (others => '0');
        P_HR_S83 <= (others => '0');
        P_HR_S84 <= (others => '0');
        P_HR_S85 <= (others => '0');
        P_HR_S86 <= (others => '0');
        P_HR_S87 <= (others => '0');
        P_HR_S88 <= (others => '0');
        P_HR_S89 <= (others => '0');
        P_HR_S90 <= (others => '0');
        P_HR_S91 <= (others => '0');
        P_HR_S92 <= (others => '0');
        P_HR_S93 <= (others => '0');
        P_HR_S94 <= (others => '0');
        P_HR_S95 <= (others => '0');
        P_HR_S96 <= (others => '0');
        P_HR_S97 <= (others => '0');
        P_HR_S98 <= (others => '0');
        P_HR_S99 <= (others => '0');
        P_HR_S100 <= (others => '0');
        P_HR_S101 <= (others => '0');
        P_HR_S102 <= (others => '0');
        P_HR_S103 <= (others => '0');
        P_HR_S104 <= (others => '0');
        P_HR_S105 <= (others => '0');
        P_HR_S106 <= (others => '0');
        P_HR_S107 <= (others => '0');
        P_HR_S108 <= (others => '0');
        P_HR_S109 <= (others => '0');
        P_HR_S110 <= (others => '0');
        P_HR_S111 <= (others => '0');
        P_HR_S112 <= (others => '0');
        P_HR_S113 <= (others => '0');
        P_HR_S114 <= (others => '0');
        P_HR_S115 <= (others => '0');
        P_HR_S116 <= (others => '0');
        P_HR_S117 <= (others => '0');
        P_HR_S118 <= (others => '0');
        P_HR_S119 <= (others => '0');
        P_HR_S120 <= (others => '0');
        P_HR_S121 <= (others => '0');
        P_HR_S122 <= (others => '0');
        P_HR_S123 <= (others => '0');
        P_HR_S124 <= (others => '0');
        P_HR_S125 <= (others => '0');
        P_HR_S126 <= (others => '0');
        P_HR_S127 <= (others => '0');
        P_HR_S128 <= (others => '0');
        P_HR_S129 <= (others => '0');
        P_HR_S130 <= (others => '0');
        P_HR_S131 <= (others => '0');
        P_HR_S132 <= (others => '0');
        P_HR_S133 <= (others => '0');
        P_HR_S134 <= (others => '0');
        P_HR_S135 <= (others => '0');
        P_HR_S136 <= (others => '0');
        P_HR_S137 <= (others => '0');
        P_HR_S138 <= (others => '0');
        P_HR_S139 <= (others => '0');
        P_HR_S140 <= (others => '0');
        P_HR_S141 <= (others => '0');
        P_HR_S142 <= (others => '0');
        P_HR_S143 <= (others => '0');
        P_HR_S144 <= (others => '0');
        P_HR_S145 <= (others => '0');
        P_HR_S146 <= (others => '0');
        P_HR_S147 <= (others => '0');
        P_HR_S148 <= (others => '0');
        P_HR_S149 <= (others => '0');
        P_HR_S150 <= (others => '0');
        P_HR_S151 <= (others => '0');
        P_HR_S152 <= (others => '0');
        P_HR_S153 <= (others => '0');
        P_HR_S154 <= (others => '0');
        P_HR_S155 <= (others => '0');
        P_HR_S156 <= (others => '0');
        P_HR_S157 <= (others => '0');
        P_HR_S158 <= (others => '0');
        P_HR_S159 <= (others => '0');
        P_HR_S160 <= (others => '0');
        P_HR_S161 <= (others => '0');
        P_HR_S162 <= (others => '0');
        P_HR_S163 <= (others => '0');
        P_HR_S164 <= (others => '0');
        P_HR_S165 <= (others => '0');
        P_HR_S166 <= (others => '0');
        P_HR_S167 <= (others => '0');
        P_HR_S168 <= (others => '0');
        P_HR_S169 <= (others => '0');
        P_HR_S170 <= (others => '0');
        P_HR_S171 <= (others => '0');
        P_HR_S172 <= (others => '0');
        P_HR_S173 <= (others => '0');
        P_HR_S174 <= (others => '0');
        P_HR_S175 <= (others => '0');
        P_HR_S176 <= (others => '0');
        P_HR_S177 <= (others => '0');
        P_HR_S178 <= (others => '0');
        P_HR_S179 <= (others => '0');
        P_HR_S180 <= (others => '0');
        P_HR_S181 <= (others => '0');
        P_HR_S182 <= (others => '0');
        P_HR_S183 <= (others => '0');
        P_HR_S184 <= (others => '0');
        P_HR_S185 <= (others => '0');
        P_HR_S186 <= (others => '0');
        P_HR_S187 <= (others => '0');
        P_HR_S188 <= (others => '0');
        P_HR_S189 <= (others => '0');
        P_HR_S190 <= (others => '0');
        P_HR_S191 <= (others => '0');
        P_HR_S192 <= (others => '0');
        P_HR_S193 <= (others => '0');
        P_HR_S194 <= (others => '0');
        P_HR_S195 <= (others => '0');
        P_HR_S196 <= (others => '0');
        P_HR_S197 <= (others => '0');
        P_HR_S198 <= (others => '0');
        P_HR_S199 <= (others => '0');
        P_HR_S200 <= (others => '0');
        P_HR_S201 <= (others => '0');
        P_HR_S202 <= (others => '0');
        P_HR_S203 <= (others => '0');
        P_HR_S204 <= (others => '0');
        P_HR_S205 <= (others => '0');
        P_HR_S206 <= (others => '0');
        P_HR_S207 <= (others => '0');
        P_HR_S208 <= (others => '0');
        P_HR_S209 <= (others => '0');
        P_HR_S210 <= (others => '0');
        P_HR_S211 <= (others => '0');
        P_HR_S212 <= (others => '0');
        P_HR_S213 <= (others => '0');
        P_HR_S214 <= (others => '0');
        P_HR_S215 <= (others => '0');
        P_HR_S216 <= (others => '0');
        P_HR_S217 <= (others => '0');
        P_HR_S218 <= (others => '0');
        P_HR_S219 <= (others => '0');
        P_HR_S220 <= (others => '0');
        P_HR_S221 <= (others => '0');
        P_HR_S222 <= (others => '0');
        P_HR_S223 <= (others => '0');
        P_HR_S224 <= (others => '0');
        P_HR_S225 <= (others => '0');
        P_HR_S226 <= (others => '0');
        P_HR_S227 <= (others => '0');
        P_HR_S228 <= (others => '0');
        P_HR_S229 <= (others => '0');
        P_HR_S230 <= (others => '0');
        P_HR_S231 <= (others => '0');
        P_HR_S232 <= (others => '0');
        P_HR_S233 <= (others => '0');
        P_HR_S234 <= (others => '0');
        P_HR_S235 <= (others => '0');
        P_HR_S236 <= (others => '0');
        P_HR_S237 <= (others => '0');
        P_HR_S238 <= (others => '0');
        P_HR_S239 <= (others => '0');
        P_HR_S240 <= (others => '0');
        P_HR_S241 <= (others => '0');
        P_HR_S242 <= (others => '0');
        P_HR_S243 <= (others => '0');
        P_HR_S244 <= (others => '0');
        P_HR_S245 <= (others => '0');
        P_HR_S246 <= (others => '0');
        P_HR_S247 <= (others => '0');
        P_HR_S248 <= (others => '0');
        P_HR_S249 <= (others => '0');
        P_HR_S250 <= (others => '0');
        P_HR_S251 <= (others => '0');
        P_HR_S252 <= (others => '0');
        P_HR_S253 <= (others => '0');
        P_HR_S254 <= (others => '0');
        P_HR_S255 <= (others => '0');
        P_HR_S256 <= (others => '0');
        P_HR_S257 <= (others => '0');
        P_HR_S258 <= (others => '0');
        P_HR_S259 <= (others => '0');
        P_HR_S260 <= (others => '0');
        P_HR_S261 <= (others => '0');
        P_HR_S262 <= (others => '0');
        P_HR_S263 <= (others => '0');
        P_HR_S264 <= (others => '0');
        P_HR_S265 <= (others => '0');
        P_HR_S266 <= (others => '0');
        P_HR_S267 <= (others => '0');
        P_HR_S268 <= (others => '0');
        P_HR_S269 <= (others => '0');
        P_HR_S270 <= (others => '0');
        P_HR_S271 <= (others => '0');
        P_HR_S272 <= (others => '0');
        P_HR_S273 <= (others => '0');
        P_HR_S274 <= (others => '0');
        P_HR_S275 <= (others => '0');
        P_HR_S276 <= (others => '0');
        P_HR_S277 <= (others => '0');
        P_HR_S278 <= (others => '0');
        P_HR_S279 <= (others => '0');
        P_HR_S280 <= (others => '0');
        P_HR_S281 <= (others => '0');
        P_HR_S282 <= (others => '0');
        P_HR_S283 <= (others => '0');
        P_HR_S284 <= (others => '0');
        P_HR_S285 <= (others => '0');
        P_HR_S286 <= (others => '0');
        P_HR_S287 <= (others => '0');
        P_HR_S288 <= (others => '0');
        P_HR_S289 <= (others => '0');
        P_HR_S290 <= (others => '0');
        P_HR_S291 <= (others => '0');
        P_HR_S292 <= (others => '0');
        P_HR_S293 <= (others => '0');
        P_HR_S294 <= (others => '0');
        P_HR_S295 <= (others => '0');
        P_HR_S296 <= (others => '0');
        P_HR_S297 <= (others => '0');
        P_HR_S298 <= (others => '0');
        P_HR_S299 <= (others => '0');
        P_HR_S300 <= (others => '0');
        P_HR_S301 <= (others => '0');
        P_HR_S302 <= (others => '0');
        P_HR_S303 <= (others => '0');
        P_HR_S304 <= (others => '0');
        P_HR_S305 <= (others => '0');
        P_HR_S306 <= (others => '0');
        P_HR_S307 <= (others => '0');
        P_HR_S308 <= (others => '0');
        P_HR_S309 <= (others => '0');
        P_HR_S310 <= (others => '0');
        P_HR_S311 <= (others => '0');
        P_HR_S312 <= (others => '0');
        P_HR_S313 <= (others => '0');
        P_HR_S314 <= (others => '0');
        P_HR_S315 <= (others => '0');
        P_HR_S316 <= (others => '0');
        P_HR_S317 <= (others => '0');
        P_HR_S318 <= (others => '0');
        P_HR_S319 <= (others => '0');
        P_HR_S320 <= (others => '0');
        P_HR_S321 <= (others => '0');
        P_HR_S322 <= (others => '0');
        P_HR_S323 <= (others => '0');
        P_HR_S324 <= (others => '0');
        P_HR_S325 <= (others => '0');
        P_HR_S326 <= (others => '0');
        P_HR_S327 <= (others => '0');
        P_HR_S328 <= (others => '0');
        P_HR_S329 <= (others => '0');
        P_HR_S330 <= (others => '0');
        P_HR_S331 <= (others => '0');
        P_HR_S332 <= (others => '0');
        P_HR_S333 <= (others => '0');
        P_HR_S334 <= (others => '0');
        P_HR_S335 <= (others => '0');
        P_HR_S336 <= (others => '0');
        P_HR_S337 <= (others => '0');
        P_HR_S338 <= (others => '0');
        P_HR_S339 <= (others => '0');
        P_HR_S340 <= (others => '0');
        P_HR_S341 <= (others => '0');
        P_HR_S342 <= (others => '0');
        P_HR_S343 <= (others => '0');
        P_HR_S344 <= (others => '0');
        P_HR_S345 <= (others => '0');
        P_HR_S346 <= (others => '0');
        P_HR_S347 <= (others => '0');
        P_HR_S348 <= (others => '0');
        P_HR_S349 <= (others => '0');
        P_HR_S350 <= (others => '0');
        P_HR_S351 <= (others => '0');
        P_HR_S352 <= (others => '0');
        P_HR_S353 <= (others => '0');
        P_HR_S354 <= (others => '0');
        P_HR_S355 <= (others => '0');
        P_HR_S356 <= (others => '0');
        P_HR_S357 <= (others => '0');
        P_HR_S358 <= (others => '0');
        P_HR_S359 <= (others => '0');
        P_HR_S360 <= (others => '0');
        P_HR_S361 <= (others => '0');
        P_HR_S362 <= (others => '0');
        P_HR_S363 <= (others => '0');
        P_HR_S364 <= (others => '0');
        P_HR_S365 <= (others => '0');
        P_HR_S366 <= (others => '0');
        P_HR_S367 <= (others => '0');
        P_HR_S368 <= (others => '0');
        P_HR_S369 <= (others => '0');
        P_HR_S370 <= (others => '0');
        P_HR_S371 <= (others => '0');
        P_HR_S372 <= (others => '0');
        P_HR_S373 <= (others => '0');
        P_HR_S374 <= (others => '0');
        P_HR_S375 <= (others => '0');
        P_HR_S376 <= (others => '0');
        P_HR_S377 <= (others => '0');
        P_HR_S378 <= (others => '0');
        P_HR_S379 <= (others => '0');
        P_HR_S380 <= (others => '0');
        P_HR_S381 <= (others => '0');
        P_HR_S382 <= (others => '0');
        P_HR_S383 <= (others => '0');
        P_HR_S384 <= (others => '0');
        P_HR_S385 <= (others => '0');
        P_HR_S386 <= (others => '0');
        P_HR_S387 <= (others => '0');
        P_HR_S388 <= (others => '0');
        P_HR_S389 <= (others => '0');
        P_HR_S390 <= (others => '0');
        P_HR_S391 <= (others => '0');
        P_HR_S392 <= (others => '0');
        P_HR_S393 <= (others => '0');
        P_HR_S394 <= (others => '0');
        P_HR_S395 <= (others => '0');
        P_HR_S396 <= (others => '0');
        P_HR_S397 <= (others => '0');
        P_HR_S398 <= (others => '0');
        P_HR_S399 <= (others => '0');
        P_HR_S400 <= (others => '0');
        P_HR_S401 <= (others => '0');
        P_HR_S402 <= (others => '0');
        P_HR_S403 <= (others => '0');
        P_HR_S404 <= (others => '0');
        P_HR_S405 <= (others => '0');
        P_HR_S406 <= (others => '0');
        P_HR_S407 <= (others => '0');
        P_HR_S408 <= (others => '0');
        P_HR_S409 <= (others => '0');
        P_HR_S410 <= (others => '0');
        P_HR_S411 <= (others => '0');
        P_HR_S412 <= (others => '0');
        P_HR_S413 <= (others => '0');
        P_HR_S414 <= (others => '0');
        P_HR_S415 <= (others => '0');
        P_HR_S416 <= (others => '0');
        P_HR_S417 <= (others => '0');
        P_HR_S418 <= (others => '0');
        P_HR_S419 <= (others => '0');
        P_HR_S420 <= (others => '0');
        P_HR_S421 <= (others => '0');
        P_HR_S422 <= (others => '0');
        P_HR_S423 <= (others => '0');
        P_HR_S424 <= (others => '0');
        P_HR_S425 <= (others => '0');
        P_HR_S426 <= (others => '0');
        P_HR_S427 <= (others => '0');
        P_HR_S428 <= (others => '0');
        P_HR_S429 <= (others => '0');
        P_HR_S430 <= (others => '0');
        P_HR_S431 <= (others => '0');
        P_HR_S432 <= (others => '0');
        P_HR_S433 <= (others => '0');
        P_HR_S434 <= (others => '0');
        P_HR_S435 <= (others => '0');
        P_HR_S436 <= (others => '0');
        P_HR_S437 <= (others => '0');
        P_HR_S438 <= (others => '0');
        P_HR_S439 <= (others => '0');
        P_HR_S440 <= (others => '0');
        P_HR_S441 <= (others => '0');
        P_HR_S442 <= (others => '0');
        P_HR_S443 <= (others => '0');
        P_HR_S444 <= (others => '0');
        P_HR_S445 <= (others => '0');
        P_HR_S446 <= (others => '0');
        P_HR_S447 <= (others => '0');
        P_HR_S448 <= (others => '0');
        P_HR_S449 <= (others => '0');
        P_HR_S450 <= (others => '0');
        P_HR_S451 <= (others => '0');
        P_HR_S452 <= (others => '0');
        P_HR_S453 <= (others => '0');
        P_HR_S454 <= (others => '0');
        P_HR_S455 <= (others => '0');
        P_HR_S456 <= (others => '0');
        P_HR_S457 <= (others => '0');
        P_HR_S458 <= (others => '0');
        P_HR_S459 <= (others => '0');
        P_HR_S460 <= (others => '0');
        P_HR_S461 <= (others => '0');
        P_HR_S462 <= (others => '0');
        P_HR_S463 <= (others => '0');
        P_HR_S464 <= (others => '0');
        P_HR_S465 <= (others => '0');
        P_HR_S466 <= (others => '0');
        P_HR_S467 <= (others => '0');
        P_HR_S468 <= (others => '0');
        P_HR_S469 <= (others => '0');
        P_HR_S470 <= (others => '0');
        P_HR_S471 <= (others => '0');
        P_HR_S472 <= (others => '0');
        P_HR_S473 <= (others => '0');
        P_HR_S474 <= (others => '0');
        P_HR_S475 <= (others => '0');
        P_HR_S476 <= (others => '0');
        P_HR_S477 <= (others => '0');
        P_HR_S478 <= (others => '0');
        P_HR_S479 <= (others => '0');
        P_HR_S480 <= (others => '0');
        P_HR_S481 <= (others => '0');
        P_HR_S482 <= (others => '0');
        P_HR_S483 <= (others => '0');
        P_HR_S484 <= (others => '0');
        P_HR_S485 <= (others => '0');
        P_HR_S486 <= (others => '0');
        P_HR_S487 <= (others => '0');
        P_HR_S488 <= (others => '0');
        P_HR_S489 <= (others => '0');
        P_HR_S490 <= (others => '0');
        P_HR_S491 <= (others => '0');
        P_HR_S492 <= (others => '0');
        P_HR_S493 <= (others => '0');
        P_HR_S494 <= (others => '0');
        P_HR_S495 <= (others => '0');
        P_HR_S496 <= (others => '0');
        P_HR_S497 <= (others => '0');
        P_HR_S498 <= (others => '0');
        P_HR_S499 <= (others => '0');
        P_HR_S500 <= (others => '0');
        P_HR_S501 <= (others => '0');
        P_HR_S502 <= (others => '0');
        P_HR_S503 <= (others => '0');
        P_HR_S504 <= (others => '0');
        P_HR_S505 <= (others => '0');
        P_HR_S506 <= (others => '0');
        P_HR_S507 <= (others => '0');
        P_HR_S508 <= (others => '0');
        P_HR_S509 <= (others => '0');
        P_HR_S510 <= (others => '0');
        P_HR_S511 <= (others => '0');
        P_HR_S512 <= (others => '0');
        P_HR_S513 <= (others => '0');
        P_HR_S514 <= (others => '0');
        P_HR_S515 <= (others => '0');
        P_HR_S516 <= (others => '0');
        P_HR_S517 <= (others => '0');
        P_HR_S518 <= (others => '0');
        P_HR_S519 <= (others => '0');
        P_HR_S520 <= (others => '0');
        P_HR_S521 <= (others => '0');
        P_HR_S522 <= (others => '0');
        P_HR_S523 <= (others => '0');
        P_HR_S524 <= (others => '0');
        P_HR_S525 <= (others => '0');
        P_HR_S526 <= (others => '0');
        P_HR_S527 <= (others => '0');
        P_HR_S528 <= (others => '0');
        P_HR_S529 <= (others => '0');
        P_HR_S530 <= (others => '0');
        P_HR_S531 <= (others => '0');
        P_HR_S532 <= (others => '0');
        P_HR_S533 <= (others => '0');
        P_HR_S534 <= (others => '0');
        P_HR_S535 <= (others => '0');
        P_HR_S536 <= (others => '0');
        P_HR_S537 <= (others => '0');
        P_HR_S538 <= (others => '0');
        P_HR_S539 <= (others => '0');
        P_HR_S540 <= (others => '0');
        P_HR_S541 <= (others => '0');
        P_HR_S542 <= (others => '0');
        P_HR_S543 <= (others => '0');
        P_HR_S544 <= (others => '0');
        P_HR_S545 <= (others => '0');
        P_HR_S546 <= (others => '0');
        P_HR_S547 <= (others => '0');
        P_HR_S548 <= (others => '0');
        P_HR_S549 <= (others => '0');
        P_HR_S550 <= (others => '0');
        P_HR_S551 <= (others => '0');
        P_HR_S552 <= (others => '0');
        P_HR_S553 <= (others => '0');
        P_HR_S554 <= (others => '0');
        P_HR_S555 <= (others => '0');
        P_HR_S556 <= (others => '0');
        P_HR_S557 <= (others => '0');
        P_HR_S558 <= (others => '0');
        P_HR_S559 <= (others => '0');
        P_HR_S560 <= (others => '0');
        P_HR_S561 <= (others => '0');
        P_HR_S562 <= (others => '0');
        P_HR_S563 <= (others => '0');
        P_HR_S564 <= (others => '0');
        P_HR_S565 <= (others => '0');
        P_HR_S566 <= (others => '0');
        P_HR_S567 <= (others => '0');
        P_HR_S568 <= (others => '0');
        P_HR_S569 <= (others => '0');
        P_HR_S570 <= (others => '0');
        P_HR_S571 <= (others => '0');
        P_HR_S572 <= (others => '0');
        P_HR_S573 <= (others => '0');
        P_HR_S574 <= (others => '0');
        P_HR_S575 <= (others => '0');
        P_HR_S576 <= (others => '0');
        P_HR_S577 <= (others => '0');
        P_HR_S578 <= (others => '0');
        P_HR_S579 <= (others => '0');
        P_HR_S580 <= (others => '0');
        P_HR_S581 <= (others => '0');
        P_HR_S582 <= (others => '0');
        P_HR_S583 <= (others => '0');
        P_HR_S584 <= (others => '0');
        P_HR_S585 <= (others => '0');
        P_HR_S586 <= (others => '0');
        P_HR_S587 <= (others => '0');
        P_HR_S588 <= (others => '0');
        P_HR_S589 <= (others => '0');
        P_HR_S590 <= (others => '0');
        P_HR_S591 <= (others => '0');
        P_HR_S592 <= (others => '0');
        P_HR_S593 <= (others => '0');
        P_HR_S594 <= (others => '0');
        P_HR_S595 <= (others => '0');
        P_HR_S596 <= (others => '0');
        P_HR_S597 <= (others => '0');
        P_HR_S598 <= (others => '0');
        P_HR_S599 <= (others => '0');
        P_HR_S600 <= (others => '0');
        P_HR_S601 <= (others => '0');
        P_HR_S602 <= (others => '0');
        P_HR_S603 <= (others => '0');
        P_HR_S604 <= (others => '0');
        P_HR_S605 <= (others => '0');
        P_HR_S606 <= (others => '0');
        P_HR_S607 <= (others => '0');
        P_HR_S608 <= (others => '0');
        P_HR_S609 <= (others => '0');
        P_HR_S610 <= (others => '0');
        P_HR_S611 <= (others => '0');
        P_HR_S612 <= (others => '0');
        P_HR_S613 <= (others => '0');
        P_HR_S614 <= (others => '0');
        P_HR_S615 <= (others => '0');
        P_HR_S616 <= (others => '0');
        P_HR_S617 <= (others => '0');
        P_HR_S618 <= (others => '0');
        P_HR_S619 <= (others => '0');
        P_HR_S620 <= (others => '0');
        P_HR_S621 <= (others => '0');
        P_HR_S622 <= (others => '0');
        P_HR_S623 <= (others => '0');
        P_HR_S624 <= (others => '0');
			
		P_TEMP_S <= (others => '0');	
		P_EDA_S <= (others => '0');	
		P_HR_S <= (others => '0');		
	    
	    stress_score <= (others => '0');
			
		elsif (rising_edge(clk)) then
		
		if (state = NORMAL) then
		
			case temp is
				when "011110111" => P_TEMP_S <= "00000000001" + P_TEMP_S1;
				when "011111000" => P_TEMP_S <= "00000111000" + P_TEMP_S2;
				when "011111001" => P_TEMP_S <= "00011010010" + P_TEMP_S3;
				when "011111010" => P_TEMP_S <= "00011000010" + P_TEMP_S4;
				when "011111011" => P_TEMP_S <= "00010011100" + P_TEMP_S5;
				when "011111100" => P_TEMP_S <= "00000000100" + P_TEMP_S6;
				when "011111101" => P_TEMP_S <= "00000000001" + P_TEMP_S7;
				when "011111110" => P_TEMP_S <= "00000111000" + P_TEMP_S8;
				when "011111111" => P_TEMP_S <= "00010011000" + P_TEMP_S9;
				when "100000000" => P_TEMP_S <= "00000111101" + P_TEMP_S10;
				when "100000001" => P_TEMP_S <= "00001000100" + P_TEMP_S11;
				when "100000010" => P_TEMP_S <= "00000101010" + P_TEMP_S12;
				when "100000011" => P_TEMP_S <= "00000010010" + P_TEMP_S13;
				when "100000100" => P_TEMP_S <= "00000001101" + P_TEMP_S14;
				when "100000101" => P_TEMP_S <= "00000001100" + P_TEMP_S15;
				when "100000110" => P_TEMP_S <= "00000001011" + P_TEMP_S16;
				when "100000111" => P_TEMP_S <= "00000001011" + P_TEMP_S17;
				when "100001000" => P_TEMP_S <= "00000001011" + P_TEMP_S18;
				when "100001001" => P_TEMP_S <= "00000100001" + P_TEMP_S19;
				when "100001010" => P_TEMP_S <= "00000101010" + P_TEMP_S20;
				when "100001011" => P_TEMP_S <= "00001000001" + P_TEMP_S21;
				when "100001100" => P_TEMP_S <= "00001001110" + P_TEMP_S22;
				when "100001101" => P_TEMP_S <= "01000111110" + P_TEMP_S23;
				when "100001110" => P_TEMP_S <= "00101001000" + P_TEMP_S24;
				when "100001111" => P_TEMP_S <= "00010100110" + P_TEMP_S25;
				when "100010000" => P_TEMP_S <= "00110010011" + P_TEMP_S26;
				when "100010001" => P_TEMP_S <= "01011111111" + P_TEMP_S27;
				when "100010010" => P_TEMP_S <= "01111111010" + P_TEMP_S28;
				when "100010011" => P_TEMP_S <= "01100000010" + P_TEMP_S29;
				when "100010100" => P_TEMP_S <= "10010010111" + P_TEMP_S30;
				when "100010101" => P_TEMP_S <= "10000111001" + P_TEMP_S31;
				when "100010110" => P_TEMP_S <= "00101100100" + P_TEMP_S32;
				when "100010111" => P_TEMP_S <= "00110101110" + P_TEMP_S33;
				when "100011000" => P_TEMP_S <= "01000010110" + P_TEMP_S34;
				when "100011001" => P_TEMP_S <= "00100101000" + P_TEMP_S35;
				when "100011010" => P_TEMP_S <= "00011101001" + P_TEMP_S36;
				when "100011011" => P_TEMP_S <= "00000110001" + P_TEMP_S37;
				when "100011100" => P_TEMP_S <= "00001111001" + P_TEMP_S38;
				when "100011101" => P_TEMP_S <= "00110010100" + P_TEMP_S39;
				when "100011110" => P_TEMP_S <= "00000000010" + P_TEMP_S40;
				when others => P_TEMP_S      <= "000000000001";
			end case;
			
			
			case eda is
				when "00001000" => P_EDA_S <= "0000000001" + P_EDA_S1;
				when "00001001" => P_EDA_S <= "0000101001" + P_EDA_S2;
				when "00001010" => P_EDA_S <= "0010010000" + P_EDA_S3;
				when "00001011" => P_EDA_S <= "0001000111" + P_EDA_S4;
				when "00001100" => P_EDA_S <= "0001100101" + P_EDA_S5;
				when "00001101" => P_EDA_S <= "0011101010" + P_EDA_S6;
				when "00001110" => P_EDA_S <= "0001110111" + P_EDA_S7;
				when "00001111" => P_EDA_S <= "0001110100" + P_EDA_S8;
				when "00010000" => P_EDA_S <= "0100100000" + P_EDA_S9;
				when "00010001" => P_EDA_S <= "0000110100" + P_EDA_S10;
				when "00010010" => P_EDA_S <= "0000010011" + P_EDA_S11;
				when "00010011" => P_EDA_S <= "0000011011" + P_EDA_S12;
				when "00010100" => P_EDA_S <= "0000011101" + P_EDA_S13;
				when "00010101" => P_EDA_S <= "0001000000" + P_EDA_S14;
				when "00010110" => P_EDA_S <= "0001011011" + P_EDA_S15;
				when "00010111" => P_EDA_S <= "0100000010" + P_EDA_S16;
				when "00011000" => P_EDA_S <= "1010001111" + P_EDA_S17;
				when "00011001" => P_EDA_S <= "0010111100" + P_EDA_S18;
				when "00011010" => P_EDA_S <= "0011000110" + P_EDA_S19;
				when "00011011" => P_EDA_S <= "0110101001" + P_EDA_S20;
				when "00011100" => P_EDA_S <= "0111000000" + P_EDA_S21;
				when "00011101" => P_EDA_S <= "0010110111" + P_EDA_S22;
				when "00011110" => P_EDA_S <= "0110011110" + P_EDA_S23;
				when "00011111" => P_EDA_S <= "0110000101" + P_EDA_S24;
				when "00100000" => P_EDA_S <= "0010011111" + P_EDA_S25;
				when "00100001" => P_EDA_S <= "0010101010" + P_EDA_S26;
				when "00100010" => P_EDA_S <= "0001100111" + P_EDA_S27;
				when "00100011" => P_EDA_S <= "0001010011" + P_EDA_S28;
				when "00100100" => P_EDA_S <= "0010000011" + P_EDA_S29;
				when "00100101" => P_EDA_S <= "0011000101" + P_EDA_S30;
				when "00100110" => P_EDA_S <= "0011010001" + P_EDA_S31;
				when "00100111" => P_EDA_S <= "0001100110" + P_EDA_S32;
				when "00101000" => P_EDA_S <= "0000110011" + P_EDA_S33;
				when "00101001" => P_EDA_S <= "0000011100" + P_EDA_S34;
				when "00101010" => P_EDA_S <= "0000010110" + P_EDA_S35;
				when "00101011" => P_EDA_S <= "0000010010" + P_EDA_S36;
				when "00101100" => P_EDA_S <= "0000010011" + P_EDA_S37;
				when "00101101" => P_EDA_S <= "0000011011" + P_EDA_S38;
				when "00101110" => P_EDA_S <= "0000011011" + P_EDA_S39;
				when "00101111" => P_EDA_S <= "0000011010" + P_EDA_S40;
				when "00110000" => P_EDA_S <= "0000011100" + P_EDA_S41;
				when "00110001" => P_EDA_S <= "0000000010" + P_EDA_S42;
				when "00110010" => P_EDA_S <= "0000000111" + P_EDA_S43;
				when "00110011" => P_EDA_S <= "0000000110" + P_EDA_S44;
				when "00110100" => P_EDA_S <= "0001100100" + P_EDA_S45;
				when "00110101" => P_EDA_S <= "0000110101" + P_EDA_S46;
				when "00110110" => P_EDA_S <= "0001100011" + P_EDA_S47;
				when "00110111" => P_EDA_S <= "0010100001" + P_EDA_S48;
				when "00111000" => P_EDA_S <= "0001100010" + P_EDA_S49;
				when "00111001" => P_EDA_S <= "0011001011" + P_EDA_S50;
				when "00111010" => P_EDA_S <= "0101100001" + P_EDA_S51;
				when "00111011" => P_EDA_S <= "0100011001" + P_EDA_S52;
				when "00111100" => P_EDA_S <= "0010000111" + P_EDA_S53;
				when "00111101" => P_EDA_S <= "0001000000" + P_EDA_S54;
				when "00111110" => P_EDA_S <= "0001000010" + P_EDA_S55;
				when "00111111" => P_EDA_S <= "0001010100" + P_EDA_S56;
				when "01000000" => P_EDA_S <= "0001001111" + P_EDA_S57;
				when "01000001" => P_EDA_S <= "0001001010" + P_EDA_S58;
				when "01000010" => P_EDA_S <= "0001000000" + P_EDA_S59;
				when "01000011" => P_EDA_S <= "0000101101" + P_EDA_S60;
				when "01000100" => P_EDA_S <= "0000110011" + P_EDA_S61;
				when "01000101" => P_EDA_S <= "0000101101" + P_EDA_S62;
				when "01000110" => P_EDA_S <= "0001001010" + P_EDA_S63;
				when "01000111" => P_EDA_S <= "0001010111" + P_EDA_S64;
				when "01001000" => P_EDA_S <= "0001010001" + P_EDA_S65;
				when "01001001" => P_EDA_S <= "0001001011" + P_EDA_S66;
				when "01001010" => P_EDA_S <= "0000110110" + P_EDA_S67;
				when "01001011" => P_EDA_S <= "0001100010" + P_EDA_S68;
				when "01001100" => P_EDA_S <= "0001101110" + P_EDA_S69;
				when "01001101" => P_EDA_S <= "0001111110" + P_EDA_S70;
				when "01001110" => P_EDA_S <= "0001011011" + P_EDA_S71;
				when "01001111" => P_EDA_S <= "0001000111" + P_EDA_S72;
				when "01010000" => P_EDA_S <= "0001000111" + P_EDA_S73;
				when "01010001" => P_EDA_S <= "0000110111" + P_EDA_S74;
				when "01010010" => P_EDA_S <= "0000110101" + P_EDA_S75;
				when "01010011" => P_EDA_S <= "0000110010" + P_EDA_S76;
				when "01010100" => P_EDA_S <= "0000111011" + P_EDA_S77;
				when "01010101" => P_EDA_S <= "0000111100" + P_EDA_S78;
				when "01010110" => P_EDA_S <= "0000011101" + P_EDA_S79;
				when "01010111" => P_EDA_S <= "0000010011" + P_EDA_S80;
				when "01011000" => P_EDA_S <= "0000001001" + P_EDA_S81;
				when "01011001" => P_EDA_S <= "0000000100" + P_EDA_S82;
				when "01011010" => P_EDA_S <= "0000000011" + P_EDA_S83;
				when "01011011" => P_EDA_S <= "0000000101" + P_EDA_S84;
				when "01011100" => P_EDA_S <= "0000000011" + P_EDA_S85;
				when "01011101" => P_EDA_S <= "0000000010" + P_EDA_S86;
				when "01011110" => P_EDA_S <= "0000000011" + P_EDA_S87;
				when "01011111" => P_EDA_S <= "0000000101" + P_EDA_S88;
				when "01100000" => P_EDA_S <= "0000000011" + P_EDA_S89;
				when "01100001" => P_EDA_S <= "0000000001" + P_EDA_S90;
				when "01111001" => P_EDA_S <= "0000000001" + P_EDA_S91;
				when "01111010" => P_EDA_S <= "0000000100" + P_EDA_S92;
				when "01111011" => P_EDA_S <= "0000000111" + P_EDA_S93;
				when "01111100" => P_EDA_S <= "0000001101" + P_EDA_S94;
				when "01111101" => P_EDA_S <= "0000011001" + P_EDA_S95;
				when "01111110" => P_EDA_S <= "0000000111" + P_EDA_S96;
				when "01111111" => P_EDA_S <= "0000001010" + P_EDA_S97;
				when "10000000" => P_EDA_S <= "0000010100" + P_EDA_S98;
				when "10000001" => P_EDA_S <= "0000001011" + P_EDA_S99;
				when "10000010" => P_EDA_S <= "0000001001" + P_EDA_S100;
				when "10000011" => P_EDA_S <= "0000001010" + P_EDA_S101;
				when "10000100" => P_EDA_S <= "0000001111" + P_EDA_S102;
				when "10000101" => P_EDA_S <= "0000100001" + P_EDA_S103;
				when "10000110" => P_EDA_S <= "0000011000" + P_EDA_S104;
				when "10000111" => P_EDA_S <= "0000011001" + P_EDA_S105;
				when "10001000" => P_EDA_S <= "0000001001" + P_EDA_S106;
				when "10001001" => P_EDA_S <= "0000000101" + P_EDA_S107;
				when "10001010" => P_EDA_S <= "0000001100" + P_EDA_S108;
				when "10001011" => P_EDA_S <= "0000001100" + P_EDA_S109;
				when "10001100" => P_EDA_S <= "0000000111" + P_EDA_S110;
				when "10001101" => P_EDA_S <= "0000010100" + P_EDA_S111;
				when "10001110" => P_EDA_S <= "0000010110" + P_EDA_S112;
				when "10001111" => P_EDA_S <= "0000010010" + P_EDA_S113;
				when "10010000" => P_EDA_S <= "0000001110" + P_EDA_S114;
				when "10010001" => P_EDA_S <= "0000010011" + P_EDA_S115;
				when "10010010" => P_EDA_S <= "0000001001" + P_EDA_S116;
				when "10010011" => P_EDA_S <= "0000011011" + P_EDA_S117;
				when "10010100" => P_EDA_S <= "0000001011" + P_EDA_S118;
				when "10010101" => P_EDA_S <= "0000001010" + P_EDA_S119;
				when "10010110" => P_EDA_S <= "0000001110" + P_EDA_S120;
				when "10010111" => P_EDA_S <= "0000001100" + P_EDA_S121;
				when "10011000" => P_EDA_S <= "0000010000" + P_EDA_S122;
				when "10011001" => P_EDA_S <= "0000001100" + P_EDA_S123;
				when "10011010" => P_EDA_S <= "0000010111" + P_EDA_S124;
				when "10011011" => P_EDA_S <= "0000010001" + P_EDA_S125;
				when "10011100" => P_EDA_S <= "0000010000" + P_EDA_S126;
				when "10011101" => P_EDA_S <= "0000001110" + P_EDA_S127;
				when "10011110" => P_EDA_S <= "0000100010" + P_EDA_S128;
				when "10011111" => P_EDA_S <= "0000111000" + P_EDA_S129;
				when "10100000" => P_EDA_S <= "0000011000" + P_EDA_S130;
				when others    => P_EDA_S <= "000000000001";
			end case;

			case hr is
				when "00000001100" => P_HR_S <= "0000001" + P_HR_S1;
				when "00000001110" => P_HR_S <= "0000001" + P_HR_S2;
				when "00000010000" => P_HR_S <= "0000010" + P_HR_S3;
				when "00000010001" => P_HR_S <= "0000001" + P_HR_S4;
				when "00000010010" => P_HR_S <= "0000001" + P_HR_S5;
				when "00000010011" => P_HR_S <= "0000001" + P_HR_S6;
				when "00000010100" => P_HR_S <= "0000001" + P_HR_S7;
				when "00000010101" => P_HR_S <= "0000001" + P_HR_S8;
				when "00000010111" => P_HR_S <= "0000001" + P_HR_S9;
				when "00000011000" => P_HR_S <= "0000001" + P_HR_S10;
				when "00000011001" => P_HR_S <= "0000001" + P_HR_S11;
				when "00000011011" => P_HR_S <= "0000001" + P_HR_S12;
				when "00000011100" => P_HR_S <= "0000001" + P_HR_S13;
				when "00000011111" => P_HR_S <= "0000010" + P_HR_S14;
				when "00000100011" => P_HR_S <= "0000001" + P_HR_S15;
				when "00000100101" => P_HR_S <= "0000001" + P_HR_S16;
				when "00000100110" => P_HR_S <= "0000001" + P_HR_S17;
				when "00000101101" => P_HR_S <= "0000001" + P_HR_S18;
				when "00000101110" => P_HR_S <= "0000010" + P_HR_S19;
				when "00000110001" => P_HR_S <= "0000001" + P_HR_S20;
				when "00000110010" => P_HR_S <= "0000001" + P_HR_S21;
				when "00000110111" => P_HR_S <= "0000001" + P_HR_S22;
				when "00000111000" => P_HR_S <= "0000010" + P_HR_S23;
				when "00000111100" => P_HR_S <= "0000001" + P_HR_S24;
				when "00001000111" => P_HR_S <= "0000001" + P_HR_S25;
				when "00001001100" => P_HR_S <= "0000001" + P_HR_S26;
				when "00001001101" => P_HR_S <= "0000001" + P_HR_S27;
				when "00001001110" => P_HR_S <= "0000001" + P_HR_S28;
				when "00001010001" => P_HR_S <= "0000001" + P_HR_S29;
				when "00001010100" => P_HR_S <= "0000001" + P_HR_S30;
				when "00001010101" => P_HR_S <= "0000010" + P_HR_S31;
				when "00001010110" => P_HR_S <= "0000001" + P_HR_S32;
				when "00001010111" => P_HR_S <= "0000001" + P_HR_S33;
				when "00001011001" => P_HR_S <= "0000010" + P_HR_S34;
				when "00001011110" => P_HR_S <= "0000001" + P_HR_S35;
				when "00001100001" => P_HR_S <= "0000001" + P_HR_S36;
				when "00001100010" => P_HR_S <= "0000001" + P_HR_S37;
				when "00001100011" => P_HR_S <= "0000001" + P_HR_S38;
				when "00001101001" => P_HR_S <= "0000001" + P_HR_S39;
				when "00001101010" => P_HR_S <= "0000001" + P_HR_S40;
				when "00001101011" => P_HR_S <= "0000001" + P_HR_S41;
				when "00001101100" => P_HR_S <= "0000010" + P_HR_S42;
				when "00001110000" => P_HR_S <= "0000001" + P_HR_S43;
				when "00001110001" => P_HR_S <= "0000001" + P_HR_S44;
				when "00001110010" => P_HR_S <= "0000001" + P_HR_S45;
				when "00001110011" => P_HR_S <= "0000001" + P_HR_S46;
				when "00001110101" => P_HR_S <= "0000001" + P_HR_S47;
				when "00001110110" => P_HR_S <= "0000010" + P_HR_S48;
				when "00001111000" => P_HR_S <= "0000001" + P_HR_S49;
				when "00001111011" => P_HR_S <= "0000001" + P_HR_S50;
				when "00001111100" => P_HR_S <= "0000001" + P_HR_S51;
				when "00001111111" => P_HR_S <= "0000011" + P_HR_S52;
				when "00010000011" => P_HR_S <= "0000001" + P_HR_S53;
				when "00010000110" => P_HR_S <= "0000001" + P_HR_S54;
				when "00010000111" => P_HR_S <= "0000001" + P_HR_S55;
				when "00010001000" => P_HR_S <= "0000001" + P_HR_S56;
				when "00010001001" => P_HR_S <= "0000001" + P_HR_S57;
				when "00010001011" => P_HR_S <= "0000001" + P_HR_S58;
				when "00010001110" => P_HR_S <= "0000001" + P_HR_S59;
				when "00010001111" => P_HR_S <= "0000011" + P_HR_S60;
				when "00010010000" => P_HR_S <= "0000011" + P_HR_S61;
				when "00010010010" => P_HR_S <= "0000001" + P_HR_S62;
				when "00010010011" => P_HR_S <= "0000001" + P_HR_S63;
				when "00010010100" => P_HR_S <= "0000001" + P_HR_S64;
				when "00010010101" => P_HR_S <= "0000001" + P_HR_S65;
				when "00010010110" => P_HR_S <= "0000001" + P_HR_S66;
				when "00010010111" => P_HR_S <= "0000010" + P_HR_S67;
				when "00010011000" => P_HR_S <= "0000001" + P_HR_S68;
				when "00010011001" => P_HR_S <= "0000001" + P_HR_S69;
				when "00010011110" => P_HR_S <= "0000001" + P_HR_S70;
				when "00010100000" => P_HR_S <= "0000001" + P_HR_S71;
				when "00010100010" => P_HR_S <= "0000001" + P_HR_S72;
				when "00010100101" => P_HR_S <= "0000001" + P_HR_S73;
				when "00010100111" => P_HR_S <= "0000001" + P_HR_S74;
				when "00010101001" => P_HR_S <= "0000001" + P_HR_S75;
				when "00010101010" => P_HR_S <= "0000010" + P_HR_S76;
				when "00010110101" => P_HR_S <= "0000001" + P_HR_S77;
				when "00010110110" => P_HR_S <= "0000010" + P_HR_S78;
				when "00010110111" => P_HR_S <= "0000001" + P_HR_S79;
				when "00010111000" => P_HR_S <= "0000001" + P_HR_S80;
				when "00010111001" => P_HR_S <= "0000001" + P_HR_S81;
				when "00010111010" => P_HR_S <= "0000001" + P_HR_S82;
				when "00010111011" => P_HR_S <= "0000010" + P_HR_S83;
				when "00010111100" => P_HR_S <= "0000001" + P_HR_S84;
				when "00010111101" => P_HR_S <= "0000001" + P_HR_S85;
				when "00010111110" => P_HR_S <= "0000001" + P_HR_S86;
				when "00010111111" => P_HR_S <= "0000001" + P_HR_S87;
				when "00011000000" => P_HR_S <= "0000010" + P_HR_S88;
				when "00011000001" => P_HR_S <= "0000001" + P_HR_S89;
				when "00011000101" => P_HR_S <= "0000010" + P_HR_S90;
				when "00011000110" => P_HR_S <= "0000011" + P_HR_S91;
				when "00011000111" => P_HR_S <= "0000001" + P_HR_S92;
				when "00011001000" => P_HR_S <= "0000001" + P_HR_S93;
				when "00011001001" => P_HR_S <= "0000001" + P_HR_S94;
				when "00011001010" => P_HR_S <= "0000011" + P_HR_S95;
				when "00011001011" => P_HR_S <= "0000010" + P_HR_S96;
				when "00011001101" => P_HR_S <= "0000011" + P_HR_S97;
				when "00011001110" => P_HR_S <= "0000010" + P_HR_S98;
				when "00011010000" => P_HR_S <= "0000010" + P_HR_S99;
				when "00011010001" => P_HR_S <= "0000010" + P_HR_S100;
				when "00011010010" => P_HR_S <= "0000001" + P_HR_S101;
				when "00011010100" => P_HR_S <= "0000001" + P_HR_S102;
				when "00011010110" => P_HR_S <= "0000001" + P_HR_S103;
				when "00011010111" => P_HR_S <= "0000001" + P_HR_S104;
				when "00011011001" => P_HR_S <= "0000001" + P_HR_S105;
				when "00011011010" => P_HR_S <= "0000001" + P_HR_S106;
				when "00011100010" => P_HR_S <= "0000001" + P_HR_S107;
				when "00011100011" => P_HR_S <= "0000001" + P_HR_S108;
				when "00011100100" => P_HR_S <= "0000001" + P_HR_S109;
				when "00011100111" => P_HR_S <= "0000001" + P_HR_S110;
				when "00011101000" => P_HR_S <= "0000001" + P_HR_S111;
				when "00011101001" => P_HR_S <= "0000001" + P_HR_S112;
				when "00011101011" => P_HR_S <= "0000001" + P_HR_S113;
				when "00011101100" => P_HR_S <= "0000001" + P_HR_S114;
				when "00011101101" => P_HR_S <= "0000001" + P_HR_S115;
				when "00011110000" => P_HR_S <= "0000001" + P_HR_S116;
				when "00011110010" => P_HR_S <= "0000001" + P_HR_S117;
				when "00011110100" => P_HR_S <= "0000001" + P_HR_S118;
				when "00011111001" => P_HR_S <= "0000001" + P_HR_S119;
				when "00011111101" => P_HR_S <= "0000001" + P_HR_S120;
				when "00100000100" => P_HR_S <= "0000001" + P_HR_S121;
				when "00100001001" => P_HR_S <= "0000001" + P_HR_S122;
				when "00100001111" => P_HR_S <= "0000001" + P_HR_S123;
				when "00100010000" => P_HR_S <= "0000011" + P_HR_S124;
				when "00100010001" => P_HR_S <= "0000001" + P_HR_S125;
				when "00100010100" => P_HR_S <= "0000001" + P_HR_S126;
				when "00100010101" => P_HR_S <= "0000001" + P_HR_S127;
				when "00100011001" => P_HR_S <= "0000001" + P_HR_S128;
				when "00100011010" => P_HR_S <= "0000001" + P_HR_S129;
				when "00100011011" => P_HR_S <= "0000001" + P_HR_S130;
				when "00100011100" => P_HR_S <= "0000001" + P_HR_S131;
				when "00100011110" => P_HR_S <= "0000001" + P_HR_S132;
				when "00100011111" => P_HR_S <= "0000001" + P_HR_S133;
				when "00100100000" => P_HR_S <= "0000100" + P_HR_S134;
				when "00100100001" => P_HR_S <= "0000001" + P_HR_S135;
				when "00100100010" => P_HR_S <= "0000001" + P_HR_S136;
				when "00100100011" => P_HR_S <= "0000001" + P_HR_S137;
				when "00100100100" => P_HR_S <= "0000001" + P_HR_S138;
				when "00100100101" => P_HR_S <= "0000001" + P_HR_S139;
				when "00100100110" => P_HR_S <= "0000001" + P_HR_S140;
				when "00100100111" => P_HR_S <= "0000001" + P_HR_S141;
				when "00100101000" => P_HR_S <= "0000011" + P_HR_S142;
				when "00100101001" => P_HR_S <= "0000001" + P_HR_S143;
				when "00100101010" => P_HR_S <= "0000011" + P_HR_S144;
				when "00100101100" => P_HR_S <= "0000010" + P_HR_S145;
				when "00100101110" => P_HR_S <= "0000001" + P_HR_S146;
				when "00100110010" => P_HR_S <= "0000001" + P_HR_S147;
				when "00100110011" => P_HR_S <= "0000001" + P_HR_S148;
				when "00100110100" => P_HR_S <= "0000001" + P_HR_S149;
				when "00100110101" => P_HR_S <= "0000001" + P_HR_S150;
				when "00100110111" => P_HR_S <= "0000010" + P_HR_S151;
				when "00100111000" => P_HR_S <= "0000001" + P_HR_S152;
				when "00100111001" => P_HR_S <= "0000011" + P_HR_S153;
				when "00100111101" => P_HR_S <= "0000011" + P_HR_S154;
				when "00101000010" => P_HR_S <= "0000001" + P_HR_S155;
				when "00101000101" => P_HR_S <= "0000001" + P_HR_S156;
				when "00101001101" => P_HR_S <= "0000001" + P_HR_S157;
				when "00101001110" => P_HR_S <= "0000001" + P_HR_S158;
				when "00101010010" => P_HR_S <= "0000001" + P_HR_S159;
				when "00101010100" => P_HR_S <= "0000001" + P_HR_S160;
				when "00101010110" => P_HR_S <= "0000001" + P_HR_S161;
				when "00101011001" => P_HR_S <= "0000001" + P_HR_S162;
				when "00101100001" => P_HR_S <= "0000001" + P_HR_S163;
				when "00101110111" => P_HR_S <= "0000001" + P_HR_S164;
				when "00110010011" => P_HR_S <= "0000001" + P_HR_S165;
				when "00110010111" => P_HR_S <= "0000001" + P_HR_S166;
				when "00110011000" => P_HR_S <= "0000001" + P_HR_S167;
				when "00110011001" => P_HR_S <= "0000001" + P_HR_S168;
				when "00110011101" => P_HR_S <= "0000001" + P_HR_S169;
				when "00110100010" => P_HR_S <= "0000001" + P_HR_S170;
				when "00110100100" => P_HR_S <= "0000001" + P_HR_S171;
				when "00110100110" => P_HR_S <= "0000010" + P_HR_S172;
				when "00110101001" => P_HR_S <= "0000001" + P_HR_S173;
				when "00110101010" => P_HR_S <= "0000001" + P_HR_S174;
				when "00110101101" => P_HR_S <= "0000001" + P_HR_S175;
				when "00110110011" => P_HR_S <= "0000011" + P_HR_S176;
				when "00110110101" => P_HR_S <= "0000001" + P_HR_S177;
				when "00110110110" => P_HR_S <= "0000011" + P_HR_S178;
				when "00110110111" => P_HR_S <= "0000001" + P_HR_S179;
				when "00110111001" => P_HR_S <= "0000001" + P_HR_S180;
				when "00110111010" => P_HR_S <= "0000001" + P_HR_S181;
				when "00110111100" => P_HR_S <= "0000011" + P_HR_S182;
				when "00110111101" => P_HR_S <= "0000001" + P_HR_S183;
				when "00110111110" => P_HR_S <= "0000001" + P_HR_S184;
				when "00111000000" => P_HR_S <= "0000001" + P_HR_S185;
				when "00111000001" => P_HR_S <= "0000010" + P_HR_S186;
				when "00111000010" => P_HR_S <= "0000001" + P_HR_S187;
				when "00111000011" => P_HR_S <= "0000001" + P_HR_S188;
				when "00111000100" => P_HR_S <= "0000010" + P_HR_S189;
				when "00111000111" => P_HR_S <= "0000011" + P_HR_S190;
				when "00111001000" => P_HR_S <= "0000001" + P_HR_S191;
				when "00111001001" => P_HR_S <= "0000010" + P_HR_S192;
				when "00111001100" => P_HR_S <= "0000001" + P_HR_S193;
				when "00111001101" => P_HR_S <= "0000001" + P_HR_S194;
				when "00111001111" => P_HR_S <= "0000011" + P_HR_S195;
				when "00111010001" => P_HR_S <= "0000001" + P_HR_S196;
				when "00111010010" => P_HR_S <= "0000001" + P_HR_S197;
				when "00111010011" => P_HR_S <= "0000010" + P_HR_S198;
				when "00111010101" => P_HR_S <= "0000001" + P_HR_S199;
				when "00111010110" => P_HR_S <= "0000001" + P_HR_S200;
				when "00111010111" => P_HR_S <= "0000011" + P_HR_S201;
				when "00111011000" => P_HR_S <= "0000001" + P_HR_S202;
				when "00111011001" => P_HR_S <= "0000011" + P_HR_S203;
				when "00111011010" => P_HR_S <= "0000001" + P_HR_S204;
				when "00111011011" => P_HR_S <= "0000001" + P_HR_S205;
				when "00111011100" => P_HR_S <= "0000011" + P_HR_S206;
				when "00111011101" => P_HR_S <= "0000100" + P_HR_S207;
				when "00111011110" => P_HR_S <= "0000010" + P_HR_S208;
				when "00111011111" => P_HR_S <= "0000011" + P_HR_S209;
				when "00111100001" => P_HR_S <= "0000011" + P_HR_S210;
				when "00111100010" => P_HR_S <= "0000001" + P_HR_S211;
				when "00111100011" => P_HR_S <= "0000001" + P_HR_S212;
				when "00111100100" => P_HR_S <= "0000001" + P_HR_S213;
				when "00111100101" => P_HR_S <= "0000010" + P_HR_S214;
				when "00111100110" => P_HR_S <= "0000100" + P_HR_S215;
				when "00111100111" => P_HR_S <= "0000010" + P_HR_S216;
				when "00111101000" => P_HR_S <= "0000001" + P_HR_S217;
				when "00111101001" => P_HR_S <= "0000010" + P_HR_S218;
				when "00111101010" => P_HR_S <= "0000010" + P_HR_S219;
				when "00111101011" => P_HR_S <= "0000001" + P_HR_S220;
				when "00111101101" => P_HR_S <= "0000110" + P_HR_S221;
				when "00111101110" => P_HR_S <= "0000001" + P_HR_S222;
				when "00111101111" => P_HR_S <= "0000011" + P_HR_S223;
				when "00111110000" => P_HR_S <= "0000011" + P_HR_S224;
				when "00111110010" => P_HR_S <= "0000011" + P_HR_S225;
				when "00111110011" => P_HR_S <= "0000011" + P_HR_S226;
				when "00111110100" => P_HR_S <= "0000001" + P_HR_S227;
				when "00111110101" => P_HR_S <= "0000010" + P_HR_S228;
				when "00111110110" => P_HR_S <= "0000110" + P_HR_S229;
				when "00111110111" => P_HR_S <= "0000010" + P_HR_S230;
				when "00111111000" => P_HR_S <= "0000110" + P_HR_S231;
				when "00111111001" => P_HR_S <= "0001010" + P_HR_S232;
				when "00111111011" => P_HR_S <= "0000001" + P_HR_S233;
				when "00111111100" => P_HR_S <= "0000111" + P_HR_S234;
				when "00111111101" => P_HR_S <= "0000010" + P_HR_S235;
				when "00111111110" => P_HR_S <= "0000001" + P_HR_S236;
				when "00111111111" => P_HR_S <= "0000011" + P_HR_S237;
				when "01000000000" => P_HR_S <= "0000001" + P_HR_S238;
				when "01000000001" => P_HR_S <= "0000001" + P_HR_S239;
				when "01000000010" => P_HR_S <= "0000001" + P_HR_S240;
				when "01000000011" => P_HR_S <= "0001000" + P_HR_S241;
				when "01000000100" => P_HR_S <= "0000011" + P_HR_S242;
				when "01000000101" => P_HR_S <= "0000001" + P_HR_S243;
				when "01000000110" => P_HR_S <= "0000010" + P_HR_S244;
				when "01000000111" => P_HR_S <= "0000110" + P_HR_S245;
				when "01000001000" => P_HR_S <= "0000011" + P_HR_S246;
				when "01000001001" => P_HR_S <= "0000011" + P_HR_S247;
				when "01000001010" => P_HR_S <= "0000001" + P_HR_S248;
				when "01000001011" => P_HR_S <= "0000111" + P_HR_S249;
				when "01000001100" => P_HR_S <= "0000011" + P_HR_S250;
				when "01000001101" => P_HR_S <= "0000110" + P_HR_S251;
				when "01000001110" => P_HR_S <= "0000001" + P_HR_S252;
				when "01000001111" => P_HR_S <= "0001111" + P_HR_S253;
				when "01000010000" => P_HR_S <= "0000110" + P_HR_S254;
				when "01000010001" => P_HR_S <= "0001100" + P_HR_S255;
				when "01000010010" => P_HR_S <= "0000111" + P_HR_S256;
				when "01000010011" => P_HR_S <= "0000010" + P_HR_S257;
				when "01000010100" => P_HR_S <= "0001110" + P_HR_S258;
				when "01000010101" => P_HR_S <= "0000101" + P_HR_S259;
				when "01000010110" => P_HR_S <= "0001000" + P_HR_S260;
				when "01000010111" => P_HR_S <= "0000111" + P_HR_S261;
				when "01000011000" => P_HR_S <= "0001001" + P_HR_S262;
				when "01000011001" => P_HR_S <= "0000110" + P_HR_S263;
				when "01000011010" => P_HR_S <= "0001010" + P_HR_S264;
				when "01000011011" => P_HR_S <= "0001000" + P_HR_S265;
				when "01000011100" => P_HR_S <= "0001000" + P_HR_S266;
				when "01000011101" => P_HR_S <= "0000110" + P_HR_S267;
				when "01000011110" => P_HR_S <= "0000101" + P_HR_S268;
				when "01000011111" => P_HR_S <= "0001000" + P_HR_S269;
				when "01000100000" => P_HR_S <= "0000110" + P_HR_S270;
				when "01000100001" => P_HR_S <= "0001001" + P_HR_S271;
				when "01000100010" => P_HR_S <= "0000110" + P_HR_S272;
				when "01000100011" => P_HR_S <= "0001001" + P_HR_S273;
				when "01000100100" => P_HR_S <= "0000100" + P_HR_S274;
				when "01000100101" => P_HR_S <= "0000011" + P_HR_S275;
				when "01000100110" => P_HR_S <= "0000101" + P_HR_S276;
				when "01000100111" => P_HR_S <= "0000011" + P_HR_S277;
				when "01000101000" => P_HR_S <= "0000111" + P_HR_S278;
				when "01000101001" => P_HR_S <= "0000110" + P_HR_S279;
				when "01000101010" => P_HR_S <= "0010101" + P_HR_S280;
				when "01000101011" => P_HR_S <= "0001011" + P_HR_S281;
				when "01000101100" => P_HR_S <= "0000111" + P_HR_S282;
				when "01000101101" => P_HR_S <= "0001100" + P_HR_S283;
				when "01000101110" => P_HR_S <= "0001100" + P_HR_S284;
				when "01000101111" => P_HR_S <= "0001100" + P_HR_S285;
				when "01000110000" => P_HR_S <= "0001001" + P_HR_S286;
				when "01000110001" => P_HR_S <= "0001001" + P_HR_S287;
				when "01000110010" => P_HR_S <= "0001001" + P_HR_S288;
				when "01000110011" => P_HR_S <= "0001010" + P_HR_S289;
				when "01000110100" => P_HR_S <= "0000100" + P_HR_S290;
				when "01000110101" => P_HR_S <= "0001100" + P_HR_S291;
				when "01000110110" => P_HR_S <= "0001011" + P_HR_S292;
				when "01000110111" => P_HR_S <= "0000110" + P_HR_S293;
				when "01000111000" => P_HR_S <= "0001000" + P_HR_S294;
				when "01000111001" => P_HR_S <= "0011101" + P_HR_S295;
				when "01000111010" => P_HR_S <= "0001110" + P_HR_S296;
				when "01000111011" => P_HR_S <= "0001100" + P_HR_S297;
				when "01000111100" => P_HR_S <= "0001010" + P_HR_S298;
				when "01000111101" => P_HR_S <= "0010001" + P_HR_S299;
				when "01000111110" => P_HR_S <= "0001100" + P_HR_S300;
				when "01000111111" => P_HR_S <= "0001000" + P_HR_S301;
				when "01001000000" => P_HR_S <= "0001000" + P_HR_S302;
				when "01001000001" => P_HR_S <= "0001100" + P_HR_S303;
				when "01001000010" => P_HR_S <= "0010000" + P_HR_S304;
				when "01001000011" => P_HR_S <= "0001011" + P_HR_S305;
				when "01001000100" => P_HR_S <= "0010001" + P_HR_S306;
				when "01001000101" => P_HR_S <= "0010000" + P_HR_S307;
				when "01001000110" => P_HR_S <= "0001011" + P_HR_S308;
				when "01001000111" => P_HR_S <= "0001001" + P_HR_S309;
				when "01001001000" => P_HR_S <= "0010000" + P_HR_S310;
				when "01001001001" => P_HR_S <= "0001001" + P_HR_S311;
				when "01001001010" => P_HR_S <= "0001100" + P_HR_S312;
				when "01001001011" => P_HR_S <= "0001010" + P_HR_S313;
				when "01001001100" => P_HR_S <= "0010011" + P_HR_S314;
				when "01001001101" => P_HR_S <= "0001100" + P_HR_S315;
				when "01001001111" => P_HR_S <= "0001110" + P_HR_S316;
				when "01001010000" => P_HR_S <= "0010011" + P_HR_S317;
				when "01001010001" => P_HR_S <= "0001001" + P_HR_S318;
				when "01001010010" => P_HR_S <= "0010011" + P_HR_S319;
				when "01001010011" => P_HR_S <= "0010101" + P_HR_S320;
				when "01001010100" => P_HR_S <= "0001111" + P_HR_S321;
				when "01001010101" => P_HR_S <= "0001011" + P_HR_S322;
				when "01001010110" => P_HR_S <= "0001101" + P_HR_S323;
				when "01001010111" => P_HR_S <= "0001111" + P_HR_S324;
				when "01001011000" => P_HR_S <= "0001101" + P_HR_S325;
				when "01001011001" => P_HR_S <= "0010001" + P_HR_S326;
				when "01001011010" => P_HR_S <= "0010011" + P_HR_S327;
				when "01001011011" => P_HR_S <= "0010000" + P_HR_S328;
				when "01001011100" => P_HR_S <= "0010000" + P_HR_S329;
				when "01001011101" => P_HR_S <= "0010110" + P_HR_S330;
				when "01001011110" => P_HR_S <= "0010110" + P_HR_S331;
				when "01001100000" => P_HR_S <= "0010011" + P_HR_S332;
				when "01001100001" => P_HR_S <= "0010001" + P_HR_S333;
				when "01001100010" => P_HR_S <= "0010110" + P_HR_S334;
				when "01001100011" => P_HR_S <= "0011001" + P_HR_S335;
				when "01001100100" => P_HR_S <= "0010011" + P_HR_S336;
				when "01001100101" => P_HR_S <= "0011001" + P_HR_S337;
				when "01001100110" => P_HR_S <= "0010010" + P_HR_S338;
				when "01001100111" => P_HR_S <= "0011000" + P_HR_S339;
				when "01001101001" => P_HR_S <= "0010010" + P_HR_S340;
				when "01001101010" => P_HR_S <= "0010110" + P_HR_S341;
				when "01001101011" => P_HR_S <= "0011010" + P_HR_S342;
				when "01001101100" => P_HR_S <= "0010010" + P_HR_S343;
				when "01001101101" => P_HR_S <= "0010110" + P_HR_S344;
				when "01001101110" => P_HR_S <= "0010101" + P_HR_S345;
				when "01001101111" => P_HR_S <= "0010110" + P_HR_S346;
				when "01001110001" => P_HR_S <= "0011010" + P_HR_S347;
				when "01001110010" => P_HR_S <= "0001101" + P_HR_S348;
				when "01001110011" => P_HR_S <= "0011000" + P_HR_S349;
				when "01001110100" => P_HR_S <= "0011000" + P_HR_S350;
				when "01001110101" => P_HR_S <= "0011100" + P_HR_S351;
				when "01001110110" => P_HR_S <= "0011010" + P_HR_S352;
				when "01001111000" => P_HR_S <= "0010001" + P_HR_S353;
				when "01001111001" => P_HR_S <= "0010011" + P_HR_S354;
				when "01001111010" => P_HR_S <= "0011010" + P_HR_S355;
				when "01001111011" => P_HR_S <= "0010110" + P_HR_S356;
				when "01001111100" => P_HR_S <= "0001111" + P_HR_S357;
				when "01001111110" => P_HR_S <= "0011000" + P_HR_S358;
				when "01001111111" => P_HR_S <= "0010001" + P_HR_S359;
				when "01010000000" => P_HR_S <= "0010001" + P_HR_S360;
				when "01010000001" => P_HR_S <= "0010100" + P_HR_S361;
				when "01010000010" => P_HR_S <= "0001000" + P_HR_S362;
				when "01010000100" => P_HR_S <= "0010000" + P_HR_S363;
				when "01010000101" => P_HR_S <= "0011001" + P_HR_S364;
				when "01010000110" => P_HR_S <= "0011111" + P_HR_S365;
				when "01010000111" => P_HR_S <= "0010101" + P_HR_S366;
				when "01010001001" => P_HR_S <= "0011110" + P_HR_S367;
				when "01010001010" => P_HR_S <= "0100100" + P_HR_S368;
				when "01010001011" => P_HR_S <= "0011001" + P_HR_S369;
				when "01010001100" => P_HR_S <= "0010101" + P_HR_S370;
				when "01010001110" => P_HR_S <= "0011010" + P_HR_S371;
				when "01010001111" => P_HR_S <= "0011111" + P_HR_S372;
				when "01010010000" => P_HR_S <= "0011000" + P_HR_S373;
				when "01010010010" => P_HR_S <= "0011101" + P_HR_S374;
				when "01010010011" => P_HR_S <= "0011010" + P_HR_S375;
				when "01010010100" => P_HR_S <= "0011010" + P_HR_S376;
				when "01010010101" => P_HR_S <= "0010011" + P_HR_S377;
				when "01010010111" => P_HR_S <= "0010101" + P_HR_S378;
				when "01010011000" => P_HR_S <= "0010111" + P_HR_S379;
				when "01010011001" => P_HR_S <= "0011110" + P_HR_S380;
				when "01010011011" => P_HR_S <= "0010111" + P_HR_S381;
				when "01010011100" => P_HR_S <= "0011011" + P_HR_S382;
				when "01010011101" => P_HR_S <= "0010111" + P_HR_S383;
				when "01010011111" => P_HR_S <= "0001111" + P_HR_S384;
				when "01010100000" => P_HR_S <= "0100001" + P_HR_S385;
				when "01010100001" => P_HR_S <= "0011110" + P_HR_S386;
				when "01010100011" => P_HR_S <= "0100111" + P_HR_S387;
				when "01010100100" => P_HR_S <= "0011011" + P_HR_S388;
				when "01010100101" => P_HR_S <= "0011010" + P_HR_S389;
				when "01010100111" => P_HR_S <= "0101000" + P_HR_S390;
				when "01010101000" => P_HR_S <= "0011001" + P_HR_S391;
				when "01010101010" => P_HR_S <= "0011011" + P_HR_S392;
				when "01010101011" => P_HR_S <= "0011100" + P_HR_S393;
				when "01010101100" => P_HR_S <= "0011111" + P_HR_S394;
				when "01010101110" => P_HR_S <= "0011011" + P_HR_S395;
				when "01010101111" => P_HR_S <= "0011110" + P_HR_S396;
				when "01010110001" => P_HR_S <= "0011100" + P_HR_S397;
				when "01010110010" => P_HR_S <= "0011100" + P_HR_S398;
				when "01010110011" => P_HR_S <= "0100001" + P_HR_S399;
				when "01010110101" => P_HR_S <= "0010001" + P_HR_S400;
				when "01010110110" => P_HR_S <= "0010101" + P_HR_S401;
				when "01010111000" => P_HR_S <= "0011101" + P_HR_S402;
				when "01010111001" => P_HR_S <= "0101000" + P_HR_S403;
				when "01010111011" => P_HR_S <= "0011101" + P_HR_S404;
				when "01010111100" => P_HR_S <= "0100011" + P_HR_S405;
				when "01010111101" => P_HR_S <= "0011111" + P_HR_S406;
				when "01010111111" => P_HR_S <= "0100000" + P_HR_S407;
				when "01011000000" => P_HR_S <= "0100011" + P_HR_S408;
				when "01011000010" => P_HR_S <= "0011110" + P_HR_S409;
				when "01011000011" => P_HR_S <= "0100011" + P_HR_S410;
				when "01011000101" => P_HR_S <= "0100001" + P_HR_S411;
				when "01011000110" => P_HR_S <= "0100001" + P_HR_S412;
				when "01011001000" => P_HR_S <= "0011100" + P_HR_S413;
				when "01011001001" => P_HR_S <= "0100001" + P_HR_S414;
				when "01011001011" => P_HR_S <= "0100011" + P_HR_S415;
				when "01011001100" => P_HR_S <= "0011111" + P_HR_S416;
				when "01011001110" => P_HR_S <= "0100001" + P_HR_S417;
				when "01011001111" => P_HR_S <= "0100101" + P_HR_S418;
				when "01011010001" => P_HR_S <= "0100011" + P_HR_S419;
				when "01011010011" => P_HR_S <= "0011111" + P_HR_S420;
				when "01011010100" => P_HR_S <= "0011111" + P_HR_S421;
				when "01011010110" => P_HR_S <= "0100011" + P_HR_S422;
				when "01011010111" => P_HR_S <= "0011011" + P_HR_S423;
				when "01011011001" => P_HR_S <= "0011100" + P_HR_S424;
				when "01011011010" => P_HR_S <= "0100101" + P_HR_S425;
				when "01011011100" => P_HR_S <= "0011010" + P_HR_S426;
				when "01011011110" => P_HR_S <= "0100100" + P_HR_S427;
				when "01011011111" => P_HR_S <= "0101010" + P_HR_S428;
				when "01011100001" => P_HR_S <= "0011111" + P_HR_S429;
				when "01011100010" => P_HR_S <= "0011111" + P_HR_S430;
				when "01011100100" => P_HR_S <= "0100011" + P_HR_S431;
				when "01011100110" => P_HR_S <= "0011111" + P_HR_S432;
				when "01011100111" => P_HR_S <= "0011111" + P_HR_S433;
				when "01011101001" => P_HR_S <= "0100001" + P_HR_S434;
				when "01011101011" => P_HR_S <= "0101001" + P_HR_S435;
				when "01011101100" => P_HR_S <= "0010111" + P_HR_S436;
				when "01011101110" => P_HR_S <= "0011000" + P_HR_S437;
				when "01011110000" => P_HR_S <= "0100011" + P_HR_S438;
				when "01011110001" => P_HR_S <= "0011101" + P_HR_S439;
				when "01011110011" => P_HR_S <= "0100000" + P_HR_S440;
				when "01011110101" => P_HR_S <= "0011001" + P_HR_S441;
				when "01011110110" => P_HR_S <= "0010110" + P_HR_S442;
				when "01011111000" => P_HR_S <= "0100001" + P_HR_S443;
				when "01011111010" => P_HR_S <= "0011010" + P_HR_S444;
				when "01011111100" => P_HR_S <= "0011100" + P_HR_S445;
				when "01011111101" => P_HR_S <= "0011111" + P_HR_S446;
				when "01011111111" => P_HR_S <= "0011001" + P_HR_S447;
				when "01100000001" => P_HR_S <= "0011100" + P_HR_S448;
				when "01100000011" => P_HR_S <= "0010111" + P_HR_S449;
				when "01100000100" => P_HR_S <= "0100001" + P_HR_S450;
				when "01100000110" => P_HR_S <= "0010100" + P_HR_S451;
				when "01100001000" => P_HR_S <= "0011010" + P_HR_S452;
				when "01100001010" => P_HR_S <= "0011001" + P_HR_S453;
				when "01100001100" => P_HR_S <= "0010101" + P_HR_S454;
				when "01100001101" => P_HR_S <= "0100100" + P_HR_S455;
				when "01100001111" => P_HR_S <= "0011000" + P_HR_S456;
				when "01100010001" => P_HR_S <= "0100100" + P_HR_S457;
				when "01100010011" => P_HR_S <= "0011111" + P_HR_S458;
				when "01100010101" => P_HR_S <= "0100001" + P_HR_S459;
				when "01100010111" => P_HR_S <= "0011010" + P_HR_S460;
				when "01100011000" => P_HR_S <= "0011100" + P_HR_S461;
				when "01100011010" => P_HR_S <= "0100011" + P_HR_S462;
				when "01100011100" => P_HR_S <= "0001100" + P_HR_S463;
				when "01100011110" => P_HR_S <= "0011111" + P_HR_S464;
				when "01100100000" => P_HR_S <= "0100000" + P_HR_S465;
				when "01100100010" => P_HR_S <= "0001101" + P_HR_S466;
				when "01100100100" => P_HR_S <= "0010100" + P_HR_S467;
				when "01100100110" => P_HR_S <= "0011011" + P_HR_S468;
				when "01100101000" => P_HR_S <= "0011010" + P_HR_S469;
				when "01100101010" => P_HR_S <= "0011010" + P_HR_S470;
				when "01100101100" => P_HR_S <= "0010111" + P_HR_S471;
				when "01100101110" => P_HR_S <= "0010110" + P_HR_S472;
				when "01100110000" => P_HR_S <= "0011010" + P_HR_S473;
				when "01100110010" => P_HR_S <= "0010110" + P_HR_S474;
				when "01100110100" => P_HR_S <= "0010100" + P_HR_S475;
				when "01100110110" => P_HR_S <= "0010110" + P_HR_S476;
				when "01100111000" => P_HR_S <= "0011100" + P_HR_S477;
				when "01100111010" => P_HR_S <= "0010101" + P_HR_S478;
				when "01100111100" => P_HR_S <= "0001101" + P_HR_S479;
				when "01100111110" => P_HR_S <= "0010001" + P_HR_S480;
				when "01101000000" => P_HR_S <= "0011001" + P_HR_S481;
				when "01101000010" => P_HR_S <= "0011000" + P_HR_S482;
				when "01101000100" => P_HR_S <= "0011000" + P_HR_S483;
				when "01101000110" => P_HR_S <= "0011000" + P_HR_S484;
				when "01101001000" => P_HR_S <= "0011000" + P_HR_S485;
				when "01101001010" => P_HR_S <= "0011011" + P_HR_S486;
				when "01101001100" => P_HR_S <= "0011000" + P_HR_S487;
				when "01101001110" => P_HR_S <= "0011001" + P_HR_S488;
				when "01101010000" => P_HR_S <= "0010110" + P_HR_S489;
				when "01101010011" => P_HR_S <= "0011110" + P_HR_S490;
				when "01101010101" => P_HR_S <= "0011000" + P_HR_S491;
				when "01101010111" => P_HR_S <= "0010001" + P_HR_S492;
				when "01101011001" => P_HR_S <= "0010011" + P_HR_S493;
				when "01101011011" => P_HR_S <= "0100010" + P_HR_S494;
				when "01101011110" => P_HR_S <= "0010110" + P_HR_S495;
				when "01101100000" => P_HR_S <= "0011100" + P_HR_S496;
				when "01101100010" => P_HR_S <= "0010110" + P_HR_S497;
				when "01101100100" => P_HR_S <= "0011010" + P_HR_S498;
				when "01101100110" => P_HR_S <= "0010111" + P_HR_S499;
				when "01101101001" => P_HR_S <= "0011100" + P_HR_S500;
				when "01101101011" => P_HR_S <= "0011001" + P_HR_S501;
				when "01101101101" => P_HR_S <= "0100001" + P_HR_S502;
				when "01101110000" => P_HR_S <= "0001111" + P_HR_S503;
				when "01101110010" => P_HR_S <= "0011100" + P_HR_S504;
				when "01101110100" => P_HR_S <= "0011111" + P_HR_S505;
				when "01101110111" => P_HR_S <= "0011000" + P_HR_S506;
				when "01101111001" => P_HR_S <= "0011100" + P_HR_S507;
				when "01101111011" => P_HR_S <= "0010011" + P_HR_S508;
				when "01101111110" => P_HR_S <= "0011011" + P_HR_S509;
				when "01110000000" => P_HR_S <= "0011000" + P_HR_S510;
				when "01110000010" => P_HR_S <= "0011001" + P_HR_S511;
				when "01110000101" => P_HR_S <= "0101011" + P_HR_S512;
				when "01110000111" => P_HR_S <= "0100101" + P_HR_S513;
				when "01110001010" => P_HR_S <= "0011100" + P_HR_S514;
				when "01110001100" => P_HR_S <= "0100011" + P_HR_S515;
				when "01110001111" => P_HR_S <= "0100001" + P_HR_S516;
				when "01110010001" => P_HR_S <= "0011100" + P_HR_S517;
				when "01110010100" => P_HR_S <= "0100010" + P_HR_S518;
				when "01110010110" => P_HR_S <= "0010001" + P_HR_S519;
				when "01110011001" => P_HR_S <= "0100011" + P_HR_S520;
				when "01110011011" => P_HR_S <= "0101011" + P_HR_S521;
				when "01110011110" => P_HR_S <= "0100010" + P_HR_S522;
				when "01110100000" => P_HR_S <= "0100101" + P_HR_S523;
				when "01110100011" => P_HR_S <= "0100101" + P_HR_S524;
				when "01110100101" => P_HR_S <= "0101010" + P_HR_S525;
				when "01110101000" => P_HR_S <= "0011000" + P_HR_S526;
				when "01110101011" => P_HR_S <= "0011111" + P_HR_S527;
				when "01110101101" => P_HR_S <= "0101001" + P_HR_S528;
				when "01110110000" => P_HR_S <= "0101111" + P_HR_S529;
				when "01110110010" => P_HR_S <= "0101110" + P_HR_S530;
				when "01110110101" => P_HR_S <= "0101101" + P_HR_S531;
				when "01110111000" => P_HR_S <= "0110001" + P_HR_S532;
				when "01110111011" => P_HR_S <= "0101010" + P_HR_S533;
				when "01110111101" => P_HR_S <= "0101001" + P_HR_S534;
				when "01111000000" => P_HR_S <= "0011111" + P_HR_S535;
				when "01111000011" => P_HR_S <= "0110000" + P_HR_S536;
				when "01111000110" => P_HR_S <= "0100001" + P_HR_S537;
				when "01111001000" => P_HR_S <= "0110101" + P_HR_S538;
				when "01111001011" => P_HR_S <= "0111100" + P_HR_S539;
				when "01111001110" => P_HR_S <= "0111100" + P_HR_S540;
				when "01111010001" => P_HR_S <= "0110011" + P_HR_S541;
				when "01111010100" => P_HR_S <= "0111010" + P_HR_S542;
				when "01111010110" => P_HR_S <= "0110011" + P_HR_S543;
				when "01111011001" => P_HR_S <= "0111111" + P_HR_S544;
				when "01111011100" => P_HR_S <= "1001100" + P_HR_S545;
				when "01111011111" => P_HR_S <= "1000000" + P_HR_S546;
				when "01111100010" => P_HR_S <= "1000111" + P_HR_S547;
				when "01111100101" => P_HR_S <= "0101001" + P_HR_S548;
				when "01111101000" => P_HR_S <= "0111100" + P_HR_S549;
				when "01111101011" => P_HR_S <= "0111110" + P_HR_S550;
				when "01111101110" => P_HR_S <= "0111000" + P_HR_S551;
				when "01111110001" => P_HR_S <= "0111100" + P_HR_S552;
				when "01111110100" => P_HR_S <= "0111010" + P_HR_S553;
				when "01111110111" => P_HR_S <= "1000000" + P_HR_S554;
				when "01111111010" => P_HR_S <= "1000000" + P_HR_S555;
				when "01111111101" => P_HR_S <= "0111010" + P_HR_S556;
				when "10000000000" => P_HR_S <= "1000011" + P_HR_S557;
				when "10000000100" => P_HR_S <= "0111000" + P_HR_S558;
				when "10000000111" => P_HR_S <= "0111010" + P_HR_S559;
				when "10000001010" => P_HR_S <= "0111000" + P_HR_S560;
				when "10000001101" => P_HR_S <= "0111101" + P_HR_S561;
				when "10000010000" => P_HR_S <= "1001010" + P_HR_S562;
				when "10000010011" => P_HR_S <= "0100001" + P_HR_S563;
				when "10000010111" => P_HR_S <= "1000011" + P_HR_S564;
				when "10000011010" => P_HR_S <= "0111011" + P_HR_S565;
				when "10000011101" => P_HR_S <= "1000101" + P_HR_S566;
				when "10000100001" => P_HR_S <= "1000000" + P_HR_S567;
				when "10000100100" => P_HR_S <= "0111101" + P_HR_S568;
				when "10000100111" => P_HR_S <= "0110001" + P_HR_S569;
				when "10000101011" => P_HR_S <= "0101011" + P_HR_S570;
				when "10000101110" => P_HR_S <= "0101110" + P_HR_S571;
				when "10000110001" => P_HR_S <= "0100111" + P_HR_S572;
				when "10000110101" => P_HR_S <= "0101010" + P_HR_S573;
				when "10000111000" => P_HR_S <= "0100011" + P_HR_S574;
				when "10000111100" => P_HR_S <= "0101010" + P_HR_S575;
				when "10000111111" => P_HR_S <= "0100100" + P_HR_S576;
				when "10001000011" => P_HR_S <= "0011011" + P_HR_S577;
				when "10001000110" => P_HR_S <= "0011010" + P_HR_S578;
				when "10001001010" => P_HR_S <= "0100011" + P_HR_S579;
				when "10001001110" => P_HR_S <= "0100011" + P_HR_S580;
				when "10001010001" => P_HR_S <= "0100111" + P_HR_S581;
				when "10001010101" => P_HR_S <= "0011100" + P_HR_S582;
				when "10001011001" => P_HR_S <= "0101011" + P_HR_S583;
				when "10001011100" => P_HR_S <= "0011011" + P_HR_S584;
				when "10001100000" => P_HR_S <= "0011101" + P_HR_S585;
				when "10001100100" => P_HR_S <= "0011011" + P_HR_S586;
				when "10001101000" => P_HR_S <= "0011111" + P_HR_S587;
				when "10001101011" => P_HR_S <= "0010100" + P_HR_S588;
				when "10001101111" => P_HR_S <= "0010110" + P_HR_S589;
				when "10001110011" => P_HR_S <= "0010001" + P_HR_S590;
				when "10001110111" => P_HR_S <= "0010011" + P_HR_S591;
				when "10001111011" => P_HR_S <= "0010001" + P_HR_S592;
				when "10001111111" => P_HR_S <= "0010111" + P_HR_S593;
				when "10010000011" => P_HR_S <= "0011000" + P_HR_S594;
				when "10010000111" => P_HR_S <= "0010000" + P_HR_S595;
				when "10010001011" => P_HR_S <= "0000110" + P_HR_S596;
				when "10010001111" => P_HR_S <= "0001111" + P_HR_S597;
				when "10010010011" => P_HR_S <= "0010001" + P_HR_S598;
				when "10010010111" => P_HR_S <= "0000101" + P_HR_S599;
				when "10010011011" => P_HR_S <= "0001001" + P_HR_S600;
				when "10010011111" => P_HR_S <= "0001000" + P_HR_S601;
				when "10010100011" => P_HR_S <= "0000011" + P_HR_S602;
				when "10010100111" => P_HR_S <= "0001000" + P_HR_S603;
				when "10010101100" => P_HR_S <= "0000110" + P_HR_S604;
				when "10010110000" => P_HR_S <= "0000110" + P_HR_S605;
				when "10010110100" => P_HR_S <= "0001011" + P_HR_S606;
				when "10010111001" => P_HR_S <= "0001000" + P_HR_S607;
				when "10010111101" => P_HR_S <= "0001000" + P_HR_S608;
				when "10011000001" => P_HR_S <= "0001100" + P_HR_S609;
				when "10011000110" => P_HR_S <= "0001100" + P_HR_S610;
				when "10011001010" => P_HR_S <= "0000110" + P_HR_S611;
				when "10011001111" => P_HR_S <= "0000110" + P_HR_S612;
				when "10011010011" => P_HR_S <= "0000011" + P_HR_S613;
				when "10011011000" => P_HR_S <= "0000011" + P_HR_S614;
				when "10011011100" => P_HR_S <= "0000101" + P_HR_S615;
				when "10011100001" => P_HR_S <= "0000010" + P_HR_S616;
				when "10011100110" => P_HR_S <= "0000010" + P_HR_S617;
				when "10011101010" => P_HR_S <= "0000001" + P_HR_S618;
				when "10011101111" => P_HR_S <= "0000001" + P_HR_S619;
				when "10100000010" => P_HR_S <= "0000001" + P_HR_S620;
				when "10100100110" => P_HR_S <= "0000001" + P_HR_S621;
				when "11001101111" => P_HR_S <= "0000001" + P_HR_S622;
				when "11010110010" => P_HR_S <= "0000001" + P_HR_S623;
				when "11011011111" => P_HR_S <= "0000001" + P_HR_S624;
				when others        => P_HR_S <= "000000000001";
			end case;
			stress_score <= P_TEMP_S * P_STRESS * P_EDA_S * P_HR_S;
		
        -- score calc
		--stress_score <= P_TEMP_S * P_STRESS * P_EDA_S * P_HR_S;
		
		elsif state = TRAINING_S then
			
			case temp is
				when "011110111" => P_TEMP_S1 <= P_TEMP_S1 + T_STRESS;
				when "011111000" => P_TEMP_S2 <= P_TEMP_S2 + T_STRESS;
				when "011111001" => P_TEMP_S3 <= P_TEMP_S3 + T_STRESS;
				when "011111010" => P_TEMP_S4 <= P_TEMP_S4 + T_STRESS;
				when "011111011" => P_TEMP_S5 <= P_TEMP_S5 + T_STRESS;
				when "011111100" => P_TEMP_S6 <= P_TEMP_S6 + T_STRESS;
				when "011111101" => P_TEMP_S7 <= P_TEMP_S7 + T_STRESS;
				when "011111110" => P_TEMP_S8 <= P_TEMP_S8 + T_STRESS;
				when "011111111" => P_TEMP_S9 <= P_TEMP_S9 + T_STRESS;
				when "100000000" => P_TEMP_S10 <= P_TEMP_S10 + T_STRESS;
				when "100000001" => P_TEMP_S11 <= P_TEMP_S11 + T_STRESS;
				when "100000010" => P_TEMP_S12 <= P_TEMP_S12 + T_STRESS;
				when "100000011" => P_TEMP_S13 <= P_TEMP_S13 + T_STRESS;
				when "100000100" => P_TEMP_S14 <= P_TEMP_S14 + T_STRESS;
				when "100000101" => P_TEMP_S15 <= P_TEMP_S15 + T_STRESS;
				when "100000110" => P_TEMP_S16 <= P_TEMP_S16 + T_STRESS;
				when "100000111" => P_TEMP_S17 <= P_TEMP_S17 + T_STRESS;
				when "100001000" => P_TEMP_S18 <= P_TEMP_S18 + T_STRESS;
				when "100001001" => P_TEMP_S19 <= P_TEMP_S19 + T_STRESS;
				when "100001010" => P_TEMP_S20 <= P_TEMP_S20 + T_STRESS;
				when "100001011" => P_TEMP_S21 <= P_TEMP_S21 + T_STRESS;
				when "100001100" => P_TEMP_S22 <= P_TEMP_S22 + T_STRESS;
				when "100001101" => P_TEMP_S23 <= P_TEMP_S23 + T_STRESS;
				when "100001110" => P_TEMP_S24 <= P_TEMP_S24 + T_STRESS;
				when "100001111" => P_TEMP_S25 <= P_TEMP_S25 + T_STRESS;
				when "100010000" => P_TEMP_S26 <= P_TEMP_S26 + T_STRESS;
				when "100010001" => P_TEMP_S27 <= P_TEMP_S27 + T_STRESS;
				when "100010010" => P_TEMP_S28 <= P_TEMP_S28 + T_STRESS;
				when "100010011" => P_TEMP_S29 <= P_TEMP_S29 + T_STRESS;
				when "100010100" => P_TEMP_S30 <= P_TEMP_S30 + T_STRESS;
				when "100010101" => P_TEMP_S31 <= P_TEMP_S31 + T_STRESS;
				when "100010110" => P_TEMP_S32 <= P_TEMP_S32 + T_STRESS;
				when "100010111" => P_TEMP_S33 <= P_TEMP_S33 + T_STRESS;
				when "100011000" => P_TEMP_S34 <= P_TEMP_S34 + T_STRESS;
				when "100011001" => P_TEMP_S35 <= P_TEMP_S35 + T_STRESS;
				when "100011010" => P_TEMP_S36 <= P_TEMP_S36 + T_STRESS;
				when "100011011" => P_TEMP_S37 <= P_TEMP_S37 + T_STRESS;
				when "100011100" => P_TEMP_S38 <= P_TEMP_S38 + T_STRESS;
				when "100011101" => P_TEMP_S39 <= P_TEMP_S39 + T_STRESS;
				when "100011110" => P_TEMP_S40 <= P_TEMP_S40 + T_STRESS;
				when  others     => null;
				
			end case;	
		
			case hr is
				when "00000001100" => P_HR_S1 <= P_HR_S1 + T_STRESS;
				when "00000001110" => P_HR_S2 <= P_HR_S2 + T_STRESS;
				when "00000010000" => P_HR_S3 <= P_HR_S3 + T_STRESS;
				when "00000010001" => P_HR_S4 <= P_HR_S4 + T_STRESS;
				when "00000010010" => P_HR_S5 <= P_HR_S5 + T_STRESS;
				when "00000010011" => P_HR_S6 <= P_HR_S6 + T_STRESS;
				when "00000010100" => P_HR_S7 <= P_HR_S7 + T_STRESS;
				when "00000010101" => P_HR_S8 <= P_HR_S8 + T_STRESS;
				when "00000010111" => P_HR_S9 <= P_HR_S9 + T_STRESS;
				when "00000011000" => P_HR_S10 <= P_HR_S10 + T_STRESS;
				when "00000011001" => P_HR_S11 <= P_HR_S11 + T_STRESS;
				when "00000011011" => P_HR_S12 <= P_HR_S12 + T_STRESS;
				when "00000011100" => P_HR_S13 <= P_HR_S13 + T_STRESS;
				when "00000011111" => P_HR_S14 <= P_HR_S14 + T_STRESS;
				when "00000100011" => P_HR_S15 <= P_HR_S15 + T_STRESS;
				when "00000100101" => P_HR_S16 <= P_HR_S16 + T_STRESS;
				when "00000100110" => P_HR_S17 <= P_HR_S17 + T_STRESS;
				when "00000101101" => P_HR_S18 <= P_HR_S18 + T_STRESS;
				when "00000101110" => P_HR_S19 <= P_HR_S19 + T_STRESS;
				when "00000110001" => P_HR_S20 <= P_HR_S20 + T_STRESS;
				when "00000110010" => P_HR_S21 <= P_HR_S21 + T_STRESS;
				when "00000110111" => P_HR_S22 <= P_HR_S22 + T_STRESS;
				when "00000111000" => P_HR_S23 <= P_HR_S23 + T_STRESS;
				when "00000111100" => P_HR_S24 <= P_HR_S24 + T_STRESS;
				when "00001000111" => P_HR_S25 <= P_HR_S25 + T_STRESS;
				when "00001001100" => P_HR_S26 <= P_HR_S26 + T_STRESS;
				when "00001001101" => P_HR_S27 <= P_HR_S27 + T_STRESS;
				when "00001001110" => P_HR_S28 <= P_HR_S28 + T_STRESS;
				when "00001010001" => P_HR_S29 <= P_HR_S29 + T_STRESS;
				when "00001010100" => P_HR_S30 <= P_HR_S30 + T_STRESS;
				when "00001010101" => P_HR_S31 <= P_HR_S31 + T_STRESS;
				when "00001010110" => P_HR_S32 <= P_HR_S32 + T_STRESS;
				when "00001010111" => P_HR_S33 <= P_HR_S33 + T_STRESS;
				when "00001011001" => P_HR_S34 <= P_HR_S34 + T_STRESS;
				when "00001011110" => P_HR_S35 <= P_HR_S35 + T_STRESS;
				when "00001100001" => P_HR_S36 <= P_HR_S36 + T_STRESS;
				when "00001100010" => P_HR_S37 <= P_HR_S37 + T_STRESS;
				when "00001100011" => P_HR_S38 <= P_HR_S38 + T_STRESS;
				when "00001101001" => P_HR_S39 <= P_HR_S39 + T_STRESS;
				when "00001101010" => P_HR_S40 <= P_HR_S40 + T_STRESS;
				when "00001101011" => P_HR_S41 <= P_HR_S41 + T_STRESS;
				when "00001101100" => P_HR_S42 <= P_HR_S42 + T_STRESS;
				when "00001110000" => P_HR_S43 <= P_HR_S43 + T_STRESS;
				when "00001110001" => P_HR_S44 <= P_HR_S44 + T_STRESS;
				when "00001110010" => P_HR_S45 <= P_HR_S45 + T_STRESS;
				when "00001110011" => P_HR_S46 <= P_HR_S46 + T_STRESS;
				when "00001110101" => P_HR_S47 <= P_HR_S47 + T_STRESS;
				when "00001110110" => P_HR_S48 <= P_HR_S48 + T_STRESS;
				when "00001111000" => P_HR_S49 <= P_HR_S49 + T_STRESS;
				when "00001111011" => P_HR_S50 <= P_HR_S50 + T_STRESS;
				when "00001111100" => P_HR_S51 <= P_HR_S51 + T_STRESS;
				when "00001111111" => P_HR_S52 <= P_HR_S52 + T_STRESS;
				when "00010000011" => P_HR_S53 <= P_HR_S53 + T_STRESS;
				when "00010000110" => P_HR_S54 <= P_HR_S54 + T_STRESS;
				when "00010000111" => P_HR_S55 <= P_HR_S55 + T_STRESS;
				when "00010001000" => P_HR_S56 <= P_HR_S56 + T_STRESS;
				when "00010001001" => P_HR_S57 <= P_HR_S57 + T_STRESS;
				when "00010001011" => P_HR_S58 <= P_HR_S58 + T_STRESS;
				when "00010001110" => P_HR_S59 <= P_HR_S59 + T_STRESS;
				when "00010001111" => P_HR_S60 <= P_HR_S60 + T_STRESS;
				when "00010010000" => P_HR_S61 <= P_HR_S61 + T_STRESS;
				when "00010010010" => P_HR_S62 <= P_HR_S62 + T_STRESS;
				when "00010010011" => P_HR_S63 <= P_HR_S63 + T_STRESS;
				when "00010010100" => P_HR_S64 <= P_HR_S64 + T_STRESS;
				when "00010010101" => P_HR_S65 <= P_HR_S65 + T_STRESS;
				when "00010010110" => P_HR_S66 <= P_HR_S66 + T_STRESS;
				when "00010010111" => P_HR_S67 <= P_HR_S67 + T_STRESS;
				when "00010011000" => P_HR_S68 <= P_HR_S68 + T_STRESS;
				when "00010011001" => P_HR_S69 <= P_HR_S69 + T_STRESS;
				when "00010011110" => P_HR_S70 <= P_HR_S70 + T_STRESS;
				when "00010100000" => P_HR_S71 <= P_HR_S71 + T_STRESS;
				when "00010100010" => P_HR_S72 <= P_HR_S72 + T_STRESS;
				when "00010100101" => P_HR_S73 <= P_HR_S73 + T_STRESS;
				when "00010100111" => P_HR_S74 <= P_HR_S74 + T_STRESS;
				when "00010101001" => P_HR_S75 <= P_HR_S75 + T_STRESS;
				when "00010101010" => P_HR_S76 <= P_HR_S76 + T_STRESS;
				when "00010110101" => P_HR_S77 <= P_HR_S77 + T_STRESS;
				when "00010110110" => P_HR_S78 <= P_HR_S78 + T_STRESS;
				when "00010110111" => P_HR_S79 <= P_HR_S79 + T_STRESS;
				when "00010111000" => P_HR_S80 <= P_HR_S80 + T_STRESS;
				when "00010111001" => P_HR_S81 <= P_HR_S81 + T_STRESS;
				when "00010111010" => P_HR_S82 <= P_HR_S82 + T_STRESS;
				when "00010111011" => P_HR_S83 <= P_HR_S83 + T_STRESS;
				when "00010111100" => P_HR_S84 <= P_HR_S84 + T_STRESS;
				when "00010111101" => P_HR_S85 <= P_HR_S85 + T_STRESS;
				when "00010111110" => P_HR_S86 <= P_HR_S86 + T_STRESS;
				when "00010111111" => P_HR_S87 <= P_HR_S87 + T_STRESS;
				when "00011000000" => P_HR_S88 <= P_HR_S88 + T_STRESS;
				when "00011000001" => P_HR_S89 <= P_HR_S89 + T_STRESS;
				when "00011000101" => P_HR_S90 <= P_HR_S90 + T_STRESS;
				when "00011000110" => P_HR_S91 <= P_HR_S91 + T_STRESS;
				when "00011000111" => P_HR_S92 <= P_HR_S92 + T_STRESS;
				when "00011001000" => P_HR_S93 <= P_HR_S93 + T_STRESS;
				when "00011001001" => P_HR_S94 <= P_HR_S94 + T_STRESS;
				when "00011001010" => P_HR_S95 <= P_HR_S95 + T_STRESS;
				when "00011001011" => P_HR_S96 <= P_HR_S96 + T_STRESS;
				when "00011001101" => P_HR_S97 <= P_HR_S97 + T_STRESS;
				when "00011001110" => P_HR_S98 <= P_HR_S98 + T_STRESS;
				when "00011010000" => P_HR_S99 <= P_HR_S99 + T_STRESS;
				when "00011010001" => P_HR_S100 <= P_HR_S100 + T_STRESS;
				when "00011010010" => P_HR_S101 <= P_HR_S101 + T_STRESS;
				when "00011010100" => P_HR_S102 <= P_HR_S102 + T_STRESS;
				when "00011010110" => P_HR_S103 <= P_HR_S103 + T_STRESS;
				when "00011010111" => P_HR_S104 <= P_HR_S104 + T_STRESS;
				when "00011011001" => P_HR_S105 <= P_HR_S105 + T_STRESS;
				when "00011011010" => P_HR_S106 <= P_HR_S106 + T_STRESS;
				when "00011100010" => P_HR_S107 <= P_HR_S107 + T_STRESS;
				when "00011100011" => P_HR_S108 <= P_HR_S108 + T_STRESS;
				when "00011100100" => P_HR_S109 <= P_HR_S109 + T_STRESS;
				when "00011100111" => P_HR_S110 <= P_HR_S110 + T_STRESS;
				when "00011101000" => P_HR_S111 <= P_HR_S111 + T_STRESS;
				when "00011101001" => P_HR_S112 <= P_HR_S112 + T_STRESS;
				when "00011101011" => P_HR_S113 <= P_HR_S113 + T_STRESS;
				when "00011101100" => P_HR_S114 <= P_HR_S114 + T_STRESS;
				when "00011101101" => P_HR_S115 <= P_HR_S115 + T_STRESS;
				when "00011110000" => P_HR_S116 <= P_HR_S116 + T_STRESS;
				when "00011110010" => P_HR_S117 <= P_HR_S117 + T_STRESS;
				when "00011110100" => P_HR_S118 <= P_HR_S118 + T_STRESS;
				when "00011111001" => P_HR_S119 <= P_HR_S119 + T_STRESS;
				when "00011111101" => P_HR_S120 <= P_HR_S120 + T_STRESS;
				when "00100000100" => P_HR_S121 <= P_HR_S121 + T_STRESS;
				when "00100001001" => P_HR_S122 <= P_HR_S122 + T_STRESS;
				when "00100001111" => P_HR_S123 <= P_HR_S123 + T_STRESS;
				when "00100010000" => P_HR_S124 <= P_HR_S124 + T_STRESS;
				when "00100010001" => P_HR_S125 <= P_HR_S125 + T_STRESS;
				when "00100010100" => P_HR_S126 <= P_HR_S126 + T_STRESS;
				when "00100010101" => P_HR_S127 <= P_HR_S127 + T_STRESS;
				when "00100011001" => P_HR_S128 <= P_HR_S128 + T_STRESS;
				when "00100011010" => P_HR_S129 <= P_HR_S129 + T_STRESS;
				when "00100011011" => P_HR_S130 <= P_HR_S130 + T_STRESS;
				when "00100011100" => P_HR_S131 <= P_HR_S131 + T_STRESS;
				when "00100011110" => P_HR_S132 <= P_HR_S132 + T_STRESS;
				when "00100011111" => P_HR_S133 <= P_HR_S133 + T_STRESS;
				when "00100100000" => P_HR_S134 <= P_HR_S134 + T_STRESS;
				when "00100100001" => P_HR_S135 <= P_HR_S135 + T_STRESS;
				when "00100100010" => P_HR_S136 <= P_HR_S136 + T_STRESS;
				when "00100100011" => P_HR_S137 <= P_HR_S137 + T_STRESS;
				when "00100100100" => P_HR_S138 <= P_HR_S138 + T_STRESS;
				when "00100100101" => P_HR_S139 <= P_HR_S139 + T_STRESS;
				when "00100100110" => P_HR_S140 <= P_HR_S140 + T_STRESS;
				when "00100100111" => P_HR_S141 <= P_HR_S141 + T_STRESS;
				when "00100101000" => P_HR_S142 <= P_HR_S142 + T_STRESS;
				when "00100101001" => P_HR_S143 <= P_HR_S143 + T_STRESS;
				when "00100101010" => P_HR_S144 <= P_HR_S144 + T_STRESS;
				when "00100101100" => P_HR_S145 <= P_HR_S145 + T_STRESS;
				when "00100101110" => P_HR_S146 <= P_HR_S146 + T_STRESS;
				when "00100110010" => P_HR_S147 <= P_HR_S147 + T_STRESS;
				when "00100110011" => P_HR_S148 <= P_HR_S148 + T_STRESS;
				when "00100110100" => P_HR_S149 <= P_HR_S149 + T_STRESS;
				when "00100110101" => P_HR_S150 <= P_HR_S150 + T_STRESS;
				when "00100110111" => P_HR_S151 <= P_HR_S151 + T_STRESS;
				when "00100111000" => P_HR_S152 <= P_HR_S152 + T_STRESS;
				when "00100111001" => P_HR_S153 <= P_HR_S153 + T_STRESS;
				when "00100111101" => P_HR_S154 <= P_HR_S154 + T_STRESS;
				when "00101000010" => P_HR_S155 <= P_HR_S155 + T_STRESS;
				when "00101000101" => P_HR_S156 <= P_HR_S156 + T_STRESS;
				when "00101001101" => P_HR_S157 <= P_HR_S157 + T_STRESS;
				when "00101001110" => P_HR_S158 <= P_HR_S158 + T_STRESS;
				when "00101010010" => P_HR_S159 <= P_HR_S159 + T_STRESS;
				when "00101010100" => P_HR_S160 <= P_HR_S160 + T_STRESS;
				when "00101010110" => P_HR_S161 <= P_HR_S161 + T_STRESS;
				when "00101011001" => P_HR_S162 <= P_HR_S162 + T_STRESS;
				when "00101100001" => P_HR_S163 <= P_HR_S163 + T_STRESS;
				when "00101110111" => P_HR_S164 <= P_HR_S164 + T_STRESS;
				when "00110010011" => P_HR_S165 <= P_HR_S165 + T_STRESS;
				when "00110010111" => P_HR_S166 <= P_HR_S166 + T_STRESS;
				when "00110011000" => P_HR_S167 <= P_HR_S167 + T_STRESS;
				when "00110011001" => P_HR_S168 <= P_HR_S168 + T_STRESS;
				when "00110011101" => P_HR_S169 <= P_HR_S169 + T_STRESS;
				when "00110100010" => P_HR_S170 <= P_HR_S170 + T_STRESS;
				when "00110100100" => P_HR_S171 <= P_HR_S171 + T_STRESS;
				when "00110100110" => P_HR_S172 <= P_HR_S172 + T_STRESS;
				when "00110101001" => P_HR_S173 <= P_HR_S173 + T_STRESS;
				when "00110101010" => P_HR_S174 <= P_HR_S174 + T_STRESS;
				when "00110101101" => P_HR_S175 <= P_HR_S175 + T_STRESS;
				when "00110110011" => P_HR_S176 <= P_HR_S176 + T_STRESS;
				when "00110110101" => P_HR_S177 <= P_HR_S177 + T_STRESS;
				when "00110110110" => P_HR_S178 <= P_HR_S178 + T_STRESS;
				when "00110110111" => P_HR_S179 <= P_HR_S179 + T_STRESS;
				when "00110111001" => P_HR_S180 <= P_HR_S180 + T_STRESS;
				when "00110111010" => P_HR_S181 <= P_HR_S181 + T_STRESS;
				when "00110111100" => P_HR_S182 <= P_HR_S182 + T_STRESS;
				when "00110111101" => P_HR_S183 <= P_HR_S183 + T_STRESS;
				when "00110111110" => P_HR_S184 <= P_HR_S184 + T_STRESS;
				when "00111000000" => P_HR_S185 <= P_HR_S185 + T_STRESS;
				when "00111000001" => P_HR_S186 <= P_HR_S186 + T_STRESS;
				when "00111000010" => P_HR_S187 <= P_HR_S187 + T_STRESS;
				when "00111000011" => P_HR_S188 <= P_HR_S188 + T_STRESS;
				when "00111000100" => P_HR_S189 <= P_HR_S189 + T_STRESS;
				when "00111000111" => P_HR_S190 <= P_HR_S190 + T_STRESS;
				when "00111001000" => P_HR_S191 <= P_HR_S191 + T_STRESS;
				when "00111001001" => P_HR_S192 <= P_HR_S192 + T_STRESS;
				when "00111001100" => P_HR_S193 <= P_HR_S193 + T_STRESS;
				when "00111001101" => P_HR_S194 <= P_HR_S194 + T_STRESS;
				when "00111001111" => P_HR_S195 <= P_HR_S195 + T_STRESS;
				when "00111010001" => P_HR_S196 <= P_HR_S196 + T_STRESS;
				when "00111010010" => P_HR_S197 <= P_HR_S197 + T_STRESS;
				when "00111010011" => P_HR_S198 <= P_HR_S198 + T_STRESS;
				when "00111010101" => P_HR_S199 <= P_HR_S199 + T_STRESS;
				when "00111010110" => P_HR_S200 <= P_HR_S200 + T_STRESS;
				when "00111010111" => P_HR_S201 <= P_HR_S201 + T_STRESS;
				when "00111011000" => P_HR_S202 <= P_HR_S202 + T_STRESS;
				when "00111011001" => P_HR_S203 <= P_HR_S203 + T_STRESS;
				when "00111011010" => P_HR_S204 <= P_HR_S204 + T_STRESS;
				when "00111011011" => P_HR_S205 <= P_HR_S205 + T_STRESS;
				when "00111011100" => P_HR_S206 <= P_HR_S206 + T_STRESS;
				when "00111011101" => P_HR_S207 <= P_HR_S207 + T_STRESS;
				when "00111011110" => P_HR_S208 <= P_HR_S208 + T_STRESS;
				when "00111011111" => P_HR_S209 <= P_HR_S209 + T_STRESS;
				when "00111100001" => P_HR_S210 <= P_HR_S210 + T_STRESS;
				when "00111100010" => P_HR_S211 <= P_HR_S211 + T_STRESS;
				when "00111100011" => P_HR_S212 <= P_HR_S212 + T_STRESS;
				when "00111100100" => P_HR_S213 <= P_HR_S213 + T_STRESS;
				when "00111100101" => P_HR_S214 <= P_HR_S214 + T_STRESS;
				when "00111100110" => P_HR_S215 <= P_HR_S215 + T_STRESS;
				when "00111100111" => P_HR_S216 <= P_HR_S216 + T_STRESS;
				when "00111101000" => P_HR_S217 <= P_HR_S217 + T_STRESS;
				when "00111101001" => P_HR_S218 <= P_HR_S218 + T_STRESS;
				when "00111101010" => P_HR_S219 <= P_HR_S219 + T_STRESS;
				when "00111101011" => P_HR_S220 <= P_HR_S220 + T_STRESS;
				when "00111101101" => P_HR_S221 <= P_HR_S221 + T_STRESS;
				when "00111101110" => P_HR_S222 <= P_HR_S222 + T_STRESS;
				when "00111101111" => P_HR_S223 <= P_HR_S223 + T_STRESS;
				when "00111110000" => P_HR_S224 <= P_HR_S224 + T_STRESS;
				when "00111110010" => P_HR_S225 <= P_HR_S225 + T_STRESS;
				when "00111110011" => P_HR_S226 <= P_HR_S226 + T_STRESS;
				when "00111110100" => P_HR_S227 <= P_HR_S227 + T_STRESS;
				when "00111110101" => P_HR_S228 <= P_HR_S228 + T_STRESS;
				when "00111110110" => P_HR_S229 <= P_HR_S229 + T_STRESS;
				when "00111110111" => P_HR_S230 <= P_HR_S230 + T_STRESS;
				when "00111111000" => P_HR_S231 <= P_HR_S231 + T_STRESS;
				when "00111111001" => P_HR_S232 <= P_HR_S232 + T_STRESS;
				when "00111111011" => P_HR_S233 <= P_HR_S233 + T_STRESS;
				when "00111111100" => P_HR_S234 <= P_HR_S234 + T_STRESS;
				when "00111111101" => P_HR_S235 <= P_HR_S235 + T_STRESS;
				when "00111111110" => P_HR_S236 <= P_HR_S236 + T_STRESS;
				when "00111111111" => P_HR_S237 <= P_HR_S237 + T_STRESS;
				when "01000000000" => P_HR_S238 <= P_HR_S238 + T_STRESS;
				when "01000000001" => P_HR_S239 <= P_HR_S239 + T_STRESS;
				when "01000000010" => P_HR_S240 <= P_HR_S240 + T_STRESS;
				when "01000000011" => P_HR_S241 <= P_HR_S241 + T_STRESS;
				when "01000000100" => P_HR_S242 <= P_HR_S242 + T_STRESS;
				when "01000000101" => P_HR_S243 <= P_HR_S243 + T_STRESS;
				when "01000000110" => P_HR_S244 <= P_HR_S244 + T_STRESS;
				when "01000000111" => P_HR_S245 <= P_HR_S245 + T_STRESS;
				when "01000001000" => P_HR_S246 <= P_HR_S246 + T_STRESS;
				when "01000001001" => P_HR_S247 <= P_HR_S247 + T_STRESS;
				when "01000001010" => P_HR_S248 <= P_HR_S248 + T_STRESS;
				when "01000001011" => P_HR_S249 <= P_HR_S249 + T_STRESS;
				when "01000001100" => P_HR_S250 <= P_HR_S250 + T_STRESS;
				when "01000001101" => P_HR_S251 <= P_HR_S251 + T_STRESS;
				when "01000001110" => P_HR_S252 <= P_HR_S252 + T_STRESS;
				when "01000001111" => P_HR_S253 <= P_HR_S253 + T_STRESS;
				when "01000010000" => P_HR_S254 <= P_HR_S254 + T_STRESS;
				when "01000010001" => P_HR_S255 <= P_HR_S255 + T_STRESS;
				when "01000010010" => P_HR_S256 <= P_HR_S256 + T_STRESS;
				when "01000010011" => P_HR_S257 <= P_HR_S257 + T_STRESS;
				when "01000010100" => P_HR_S258 <= P_HR_S258 + T_STRESS;
				when "01000010101" => P_HR_S259 <= P_HR_S259 + T_STRESS;
				when "01000010110" => P_HR_S260 <= P_HR_S260 + T_STRESS;
				when "01000010111" => P_HR_S261 <= P_HR_S261 + T_STRESS;
				when "01000011000" => P_HR_S262 <= P_HR_S262 + T_STRESS;
				when "01000011001" => P_HR_S263 <= P_HR_S263 + T_STRESS;
				when "01000011010" => P_HR_S264 <= P_HR_S264 + T_STRESS;
				when "01000011011" => P_HR_S265 <= P_HR_S265 + T_STRESS;
				when "01000011100" => P_HR_S266 <= P_HR_S266 + T_STRESS;
				when "01000011101" => P_HR_S267 <= P_HR_S267 + T_STRESS;
				when "01000011110" => P_HR_S268 <= P_HR_S268 + T_STRESS;
				when "01000011111" => P_HR_S269 <= P_HR_S269 + T_STRESS;
				when "01000100000" => P_HR_S270 <= P_HR_S270 + T_STRESS;
				when "01000100001" => P_HR_S271 <= P_HR_S271 + T_STRESS;
				when "01000100010" => P_HR_S272 <= P_HR_S272 + T_STRESS;
				when "01000100011" => P_HR_S273 <= P_HR_S273 + T_STRESS;
				when "01000100100" => P_HR_S274 <= P_HR_S274 + T_STRESS;
				when "01000100101" => P_HR_S275 <= P_HR_S275 + T_STRESS;
				when "01000100110" => P_HR_S276 <= P_HR_S276 + T_STRESS;
				when "01000100111" => P_HR_S277 <= P_HR_S277 + T_STRESS;
				when "01000101000" => P_HR_S278 <= P_HR_S278 + T_STRESS;
				when "01000101001" => P_HR_S279 <= P_HR_S279 + T_STRESS;
				when "01000101010" => P_HR_S280 <= P_HR_S280 + T_STRESS;
				when "01000101011" => P_HR_S281 <= P_HR_S281 + T_STRESS;
				when "01000101100" => P_HR_S282 <= P_HR_S282 + T_STRESS;
				when "01000101101" => P_HR_S283 <= P_HR_S283 + T_STRESS;
				when "01000101110" => P_HR_S284 <= P_HR_S284 + T_STRESS;
				when "01000101111" => P_HR_S285 <= P_HR_S285 + T_STRESS;
				when "01000110000" => P_HR_S286 <= P_HR_S286 + T_STRESS;
				when "01000110001" => P_HR_S287 <= P_HR_S287 + T_STRESS;
				when "01000110010" => P_HR_S288 <= P_HR_S288 + T_STRESS;
				when "01000110011" => P_HR_S289 <= P_HR_S289 + T_STRESS;
				when "01000110100" => P_HR_S290 <= P_HR_S290 + T_STRESS;
				when "01000110101" => P_HR_S291 <= P_HR_S291 + T_STRESS;
				when "01000110110" => P_HR_S292 <= P_HR_S292 + T_STRESS;
				when "01000110111" => P_HR_S293 <= P_HR_S293 + T_STRESS;
				when "01000111000" => P_HR_S294 <= P_HR_S294 + T_STRESS;
				when "01000111001" => P_HR_S295 <= P_HR_S295 + T_STRESS;
				when "01000111010" => P_HR_S296 <= P_HR_S296 + T_STRESS;
				when "01000111011" => P_HR_S297 <= P_HR_S297 + T_STRESS;
				when "01000111100" => P_HR_S298 <= P_HR_S298 + T_STRESS;
				when "01000111101" => P_HR_S299 <= P_HR_S299 + T_STRESS;
				when "01000111110" => P_HR_S300 <= P_HR_S300 + T_STRESS;
				when "01000111111" => P_HR_S301 <= P_HR_S301 + T_STRESS;
				when "01001000000" => P_HR_S302 <= P_HR_S302 + T_STRESS;
				when "01001000001" => P_HR_S303 <= P_HR_S303 + T_STRESS;
				when "01001000010" => P_HR_S304 <= P_HR_S304 + T_STRESS;
				when "01001000011" => P_HR_S305 <= P_HR_S305 + T_STRESS;
				when "01001000100" => P_HR_S306 <= P_HR_S306 + T_STRESS;
				when "01001000101" => P_HR_S307 <= P_HR_S307 + T_STRESS;
				when "01001000110" => P_HR_S308 <= P_HR_S308 + T_STRESS;
				when "01001000111" => P_HR_S309 <= P_HR_S309 + T_STRESS;
				when "01001001000" => P_HR_S310 <= P_HR_S310 + T_STRESS;
				when "01001001001" => P_HR_S311 <= P_HR_S311 + T_STRESS;
				when "01001001010" => P_HR_S312 <= P_HR_S312 + T_STRESS;
				when "01001001011" => P_HR_S313 <= P_HR_S313 + T_STRESS;
				when "01001001100" => P_HR_S314 <= P_HR_S314 + T_STRESS;
				when "01001001101" => P_HR_S315 <= P_HR_S315 + T_STRESS;
				when "01001001111" => P_HR_S316 <= P_HR_S316 + T_STRESS;
				when "01001010000" => P_HR_S317 <= P_HR_S317 + T_STRESS;
				when "01001010001" => P_HR_S318 <= P_HR_S318 + T_STRESS;
				when "01001010010" => P_HR_S319 <= P_HR_S319 + T_STRESS;
				when "01001010011" => P_HR_S320 <= P_HR_S320 + T_STRESS;
				when "01001010100" => P_HR_S321 <= P_HR_S321 + T_STRESS;
				when "01001010101" => P_HR_S322 <= P_HR_S322 + T_STRESS;
				when "01001010110" => P_HR_S323 <= P_HR_S323 + T_STRESS;
				when "01001010111" => P_HR_S324 <= P_HR_S324 + T_STRESS;
				when "01001011000" => P_HR_S325 <= P_HR_S325 + T_STRESS;
				when "01001011001" => P_HR_S326 <= P_HR_S326 + T_STRESS;
				when "01001011010" => P_HR_S327 <= P_HR_S327 + T_STRESS;
				when "01001011011" => P_HR_S328 <= P_HR_S328 + T_STRESS;
				when "01001011100" => P_HR_S329 <= P_HR_S329 + T_STRESS;
				when "01001011101" => P_HR_S330 <= P_HR_S330 + T_STRESS;
				when "01001011110" => P_HR_S331 <= P_HR_S331 + T_STRESS;
				when "01001100000" => P_HR_S332 <= P_HR_S332 + T_STRESS;
				when "01001100001" => P_HR_S333 <= P_HR_S333 + T_STRESS;
				when "01001100010" => P_HR_S334 <= P_HR_S334 + T_STRESS;
				when "01001100011" => P_HR_S335 <= P_HR_S335 + T_STRESS;
				when "01001100100" => P_HR_S336 <= P_HR_S336 + T_STRESS;
				when "01001100101" => P_HR_S337 <= P_HR_S337 + T_STRESS;
				when "01001100110" => P_HR_S338 <= P_HR_S338 + T_STRESS;
				when "01001100111" => P_HR_S339 <= P_HR_S339 + T_STRESS;
				when "01001101001" => P_HR_S340 <= P_HR_S340 + T_STRESS;
				when "01001101010" => P_HR_S341 <= P_HR_S341 + T_STRESS;
				when "01001101011" => P_HR_S342 <= P_HR_S342 + T_STRESS;
				when "01001101100" => P_HR_S343 <= P_HR_S343 + T_STRESS;
				when "01001101101" => P_HR_S344 <= P_HR_S344 + T_STRESS;
				when "01001101110" => P_HR_S345 <= P_HR_S345 + T_STRESS;
				when "01001101111" => P_HR_S346 <= P_HR_S346 + T_STRESS;
				when "01001110001" => P_HR_S347 <= P_HR_S347 + T_STRESS;
				when "01001110010" => P_HR_S348 <= P_HR_S348 + T_STRESS;
				when "01001110011" => P_HR_S349 <= P_HR_S349 + T_STRESS;
				when "01001110100" => P_HR_S350 <= P_HR_S350 + T_STRESS;
				when "01001110101" => P_HR_S351 <= P_HR_S351 + T_STRESS;
				when "01001110110" => P_HR_S352 <= P_HR_S352 + T_STRESS;
				when "01001111000" => P_HR_S353 <= P_HR_S353 + T_STRESS;
				when "01001111001" => P_HR_S354 <= P_HR_S354 + T_STRESS;
				when "01001111010" => P_HR_S355 <= P_HR_S355 + T_STRESS;
				when "01001111011" => P_HR_S356 <= P_HR_S356 + T_STRESS;
				when "01001111100" => P_HR_S357 <= P_HR_S357 + T_STRESS;
				when "01001111110" => P_HR_S358 <= P_HR_S358 + T_STRESS;
				when "01001111111" => P_HR_S359 <= P_HR_S359 + T_STRESS;
				when "01010000000" => P_HR_S360 <= P_HR_S360 + T_STRESS;
				when "01010000001" => P_HR_S361 <= P_HR_S361 + T_STRESS;
				when "01010000010" => P_HR_S362 <= P_HR_S362 + T_STRESS;
				when "01010000100" => P_HR_S363 <= P_HR_S363 + T_STRESS;
				when "01010000101" => P_HR_S364 <= P_HR_S364 + T_STRESS;
				when "01010000110" => P_HR_S365 <= P_HR_S365 + T_STRESS;
				when "01010000111" => P_HR_S366 <= P_HR_S366 + T_STRESS;
				when "01010001001" => P_HR_S367 <= P_HR_S367 + T_STRESS;
				when "01010001010" => P_HR_S368 <= P_HR_S368 + T_STRESS;
				when "01010001011" => P_HR_S369 <= P_HR_S369 + T_STRESS;
				when "01010001100" => P_HR_S370 <= P_HR_S370 + T_STRESS;
				when "01010001110" => P_HR_S371 <= P_HR_S371 + T_STRESS;
				when "01010001111" => P_HR_S372 <= P_HR_S372 + T_STRESS;
				when "01010010000" => P_HR_S373 <= P_HR_S373 + T_STRESS;
				when "01010010010" => P_HR_S374 <= P_HR_S374 + T_STRESS;
				when "01010010011" => P_HR_S375 <= P_HR_S375 + T_STRESS;
				when "01010010100" => P_HR_S376 <= P_HR_S376 + T_STRESS;
				when "01010010101" => P_HR_S377 <= P_HR_S377 + T_STRESS;
				when "01010010111" => P_HR_S378 <= P_HR_S378 + T_STRESS;
				when "01010011000" => P_HR_S379 <= P_HR_S379 + T_STRESS;
				when "01010011001" => P_HR_S380 <= P_HR_S380 + T_STRESS;
				when "01010011011" => P_HR_S381 <= P_HR_S381 + T_STRESS;
				when "01010011100" => P_HR_S382 <= P_HR_S382 + T_STRESS;
				when "01010011101" => P_HR_S383 <= P_HR_S383 + T_STRESS;
				when "01010011111" => P_HR_S384 <= P_HR_S384 + T_STRESS;
				when "01010100000" => P_HR_S385 <= P_HR_S385 + T_STRESS;
				when "01010100001" => P_HR_S386 <= P_HR_S386 + T_STRESS;
				when "01010100011" => P_HR_S387 <= P_HR_S387 + T_STRESS;
				when "01010100100" => P_HR_S388 <= P_HR_S388 + T_STRESS;
				when "01010100101" => P_HR_S389 <= P_HR_S389 + T_STRESS;
				when "01010100111" => P_HR_S390 <= P_HR_S390 + T_STRESS;
				when "01010101000" => P_HR_S391 <= P_HR_S391 + T_STRESS;
				when "01010101010" => P_HR_S392 <= P_HR_S392 + T_STRESS;
				when "01010101011" => P_HR_S393 <= P_HR_S393 + T_STRESS;
				when "01010101100" => P_HR_S394 <= P_HR_S394 + T_STRESS;
				when "01010101110" => P_HR_S395 <= P_HR_S395 + T_STRESS;
				when "01010101111" => P_HR_S396 <= P_HR_S396 + T_STRESS;
				when "01010110001" => P_HR_S397 <= P_HR_S397 + T_STRESS;
				when "01010110010" => P_HR_S398 <= P_HR_S398 + T_STRESS;
				when "01010110011" => P_HR_S399 <= P_HR_S399 + T_STRESS;
				when "01010110101" => P_HR_S400 <= P_HR_S400 + T_STRESS;
				when "01010110110" => P_HR_S401 <= P_HR_S401 + T_STRESS;
				when "01010111000" => P_HR_S402 <= P_HR_S402 + T_STRESS;
				when "01010111001" => P_HR_S403 <= P_HR_S403 + T_STRESS;
				when "01010111011" => P_HR_S404 <= P_HR_S404 + T_STRESS;
				when "01010111100" => P_HR_S405 <= P_HR_S405 + T_STRESS;
				when "01010111101" => P_HR_S406 <= P_HR_S406 + T_STRESS;
				when "01010111111" => P_HR_S407 <= P_HR_S407 + T_STRESS;
				when "01011000000" => P_HR_S408 <= P_HR_S408 + T_STRESS;
				when "01011000010" => P_HR_S409 <= P_HR_S409 + T_STRESS;
				when "01011000011" => P_HR_S410 <= P_HR_S410 + T_STRESS;
				when "01011000101" => P_HR_S411 <= P_HR_S411 + T_STRESS;
				when "01011000110" => P_HR_S412 <= P_HR_S412 + T_STRESS;
				when "01011001000" => P_HR_S413 <= P_HR_S413 + T_STRESS;
				when "01011001001" => P_HR_S414 <= P_HR_S414 + T_STRESS;
				when "01011001011" => P_HR_S415 <= P_HR_S415 + T_STRESS;
				when "01011001100" => P_HR_S416 <= P_HR_S416 + T_STRESS;
				when "01011001110" => P_HR_S417 <= P_HR_S417 + T_STRESS;
				when "01011001111" => P_HR_S418 <= P_HR_S418 + T_STRESS;
				when "01011010001" => P_HR_S419 <= P_HR_S419 + T_STRESS;
				when "01011010011" => P_HR_S420 <= P_HR_S420 + T_STRESS;
				when "01011010100" => P_HR_S421 <= P_HR_S421 + T_STRESS;
				when "01011010110" => P_HR_S422 <= P_HR_S422 + T_STRESS;
				when "01011010111" => P_HR_S423 <= P_HR_S423 + T_STRESS;
				when "01011011001" => P_HR_S424 <= P_HR_S424 + T_STRESS;
				when "01011011010" => P_HR_S425 <= P_HR_S425 + T_STRESS;
				when "01011011100" => P_HR_S426 <= P_HR_S426 + T_STRESS;
				when "01011011110" => P_HR_S427 <= P_HR_S427 + T_STRESS;
				when "01011011111" => P_HR_S428 <= P_HR_S428 + T_STRESS;
				when "01011100001" => P_HR_S429 <= P_HR_S429 + T_STRESS;
				when "01011100010" => P_HR_S430 <= P_HR_S430 + T_STRESS;
				when "01011100100" => P_HR_S431 <= P_HR_S431 + T_STRESS;
				when "01011100110" => P_HR_S432 <= P_HR_S432 + T_STRESS;
				when "01011100111" => P_HR_S433 <= P_HR_S433 + T_STRESS;
				when "01011101001" => P_HR_S434 <= P_HR_S434 + T_STRESS;
				when "01011101011" => P_HR_S435 <= P_HR_S435 + T_STRESS;
				when "01011101100" => P_HR_S436 <= P_HR_S436 + T_STRESS;
				when "01011101110" => P_HR_S437 <= P_HR_S437 + T_STRESS;
				when "01011110000" => P_HR_S438 <= P_HR_S438 + T_STRESS;
				when "01011110001" => P_HR_S439 <= P_HR_S439 + T_STRESS;
				when "01011110011" => P_HR_S440 <= P_HR_S440 + T_STRESS;
				when "01011110101" => P_HR_S441 <= P_HR_S441 + T_STRESS;
				when "01011110110" => P_HR_S442 <= P_HR_S442 + T_STRESS;
				when "01011111000" => P_HR_S443 <= P_HR_S443 + T_STRESS;
				when "01011111010" => P_HR_S444 <= P_HR_S444 + T_STRESS;
				when "01011111100" => P_HR_S445 <= P_HR_S445 + T_STRESS;
				when "01011111101" => P_HR_S446 <= P_HR_S446 + T_STRESS;
				when "01011111111" => P_HR_S447 <= P_HR_S447 + T_STRESS;
				when "01100000001" => P_HR_S448 <= P_HR_S448 + T_STRESS;
				when "01100000011" => P_HR_S449 <= P_HR_S449 + T_STRESS;
				when "01100000100" => P_HR_S450 <= P_HR_S450 + T_STRESS;
				when "01100000110" => P_HR_S451 <= P_HR_S451 + T_STRESS;
				when "01100001000" => P_HR_S452 <= P_HR_S452 + T_STRESS;
				when "01100001010" => P_HR_S453 <= P_HR_S453 + T_STRESS;
				when "01100001100" => P_HR_S454 <= P_HR_S454 + T_STRESS;
				when "01100001101" => P_HR_S455 <= P_HR_S455 + T_STRESS;
				when "01100001111" => P_HR_S456 <= P_HR_S456 + T_STRESS;
				when "01100010001" => P_HR_S457 <= P_HR_S457 + T_STRESS;
				when "01100010011" => P_HR_S458 <= P_HR_S458 + T_STRESS;
				when "01100010101" => P_HR_S459 <= P_HR_S459 + T_STRESS;
				when "01100010111" => P_HR_S460 <= P_HR_S460 + T_STRESS;
				when "01100011000" => P_HR_S461 <= P_HR_S461 + T_STRESS;
				when "01100011010" => P_HR_S462 <= P_HR_S462 + T_STRESS;
				when "01100011100" => P_HR_S463 <= P_HR_S463 + T_STRESS;
				when "01100011110" => P_HR_S464 <= P_HR_S464 + T_STRESS;
				when "01100100000" => P_HR_S465 <= P_HR_S465 + T_STRESS;
				when "01100100010" => P_HR_S466 <= P_HR_S466 + T_STRESS;
				when "01100100100" => P_HR_S467 <= P_HR_S467 + T_STRESS;
				when "01100100110" => P_HR_S468 <= P_HR_S468 + T_STRESS;
				when "01100101000" => P_HR_S469 <= P_HR_S469 + T_STRESS;
				when "01100101010" => P_HR_S470 <= P_HR_S470 + T_STRESS;
				when "01100101100" => P_HR_S471 <= P_HR_S471 + T_STRESS;
				when "01100101110" => P_HR_S472 <= P_HR_S472 + T_STRESS;
				when "01100110000" => P_HR_S473 <= P_HR_S473 + T_STRESS;
				when "01100110010" => P_HR_S474 <= P_HR_S474 + T_STRESS;
				when "01100110100" => P_HR_S475 <= P_HR_S475 + T_STRESS;
				when "01100110110" => P_HR_S476 <= P_HR_S476 + T_STRESS;
				when "01100111000" => P_HR_S477 <= P_HR_S477 + T_STRESS;
				when "01100111010" => P_HR_S478 <= P_HR_S478 + T_STRESS;
				when "01100111100" => P_HR_S479 <= P_HR_S479 + T_STRESS;
				when "01100111110" => P_HR_S480 <= P_HR_S480 + T_STRESS;
				when "01101000000" => P_HR_S481 <= P_HR_S481 + T_STRESS;
				when "01101000010" => P_HR_S482 <= P_HR_S482 + T_STRESS;
				when "01101000100" => P_HR_S483 <= P_HR_S483 + T_STRESS;
				when "01101000110" => P_HR_S484 <= P_HR_S484 + T_STRESS;
				when "01101001000" => P_HR_S485 <= P_HR_S485 + T_STRESS;
				when "01101001010" => P_HR_S486 <= P_HR_S486 + T_STRESS;
				when "01101001100" => P_HR_S487 <= P_HR_S487 + T_STRESS;
				when "01101001110" => P_HR_S488 <= P_HR_S488 + T_STRESS;
				when "01101010000" => P_HR_S489 <= P_HR_S489 + T_STRESS;
				when "01101010011" => P_HR_S490 <= P_HR_S490 + T_STRESS;
				when "01101010101" => P_HR_S491 <= P_HR_S491 + T_STRESS;
				when "01101010111" => P_HR_S492 <= P_HR_S492 + T_STRESS;
				when "01101011001" => P_HR_S493 <= P_HR_S493 + T_STRESS;
				when "01101011011" => P_HR_S494 <= P_HR_S494 + T_STRESS;
				when "01101011110" => P_HR_S495 <= P_HR_S495 + T_STRESS;
				when "01101100000" => P_HR_S496 <= P_HR_S496 + T_STRESS;
				when "01101100010" => P_HR_S497 <= P_HR_S497 + T_STRESS;
				when "01101100100" => P_HR_S498 <= P_HR_S498 + T_STRESS;
				when "01101100110" => P_HR_S499 <= P_HR_S499 + T_STRESS;
				when "01101101001" => P_HR_S500 <= P_HR_S500 + T_STRESS;
				when "01101101011" => P_HR_S501 <= P_HR_S501 + T_STRESS;
				when "01101101101" => P_HR_S502 <= P_HR_S502 + T_STRESS;
				when "01101110000" => P_HR_S503 <= P_HR_S503 + T_STRESS;
				when "01101110010" => P_HR_S504 <= P_HR_S504 + T_STRESS;
				when "01101110100" => P_HR_S505 <= P_HR_S505 + T_STRESS;
				when "01101110111" => P_HR_S506 <= P_HR_S506 + T_STRESS;
				when "01101111001" => P_HR_S507 <= P_HR_S507 + T_STRESS;
				when "01101111011" => P_HR_S508 <= P_HR_S508 + T_STRESS;
				when "01101111110" => P_HR_S509 <= P_HR_S509 + T_STRESS;
				when "01110000000" => P_HR_S510 <= P_HR_S510 + T_STRESS;
				when "01110000010" => P_HR_S511 <= P_HR_S511 + T_STRESS;
				when "01110000101" => P_HR_S512 <= P_HR_S512 + T_STRESS;
				when "01110000111" => P_HR_S513 <= P_HR_S513 + T_STRESS;
				when "01110001010" => P_HR_S514 <= P_HR_S514 + T_STRESS;
				when "01110001100" => P_HR_S515 <= P_HR_S515 + T_STRESS;
				when "01110001111" => P_HR_S516 <= P_HR_S516 + T_STRESS;
				when "01110010001" => P_HR_S517 <= P_HR_S517 + T_STRESS;
				when "01110010100" => P_HR_S518 <= P_HR_S518 + T_STRESS;
				when "01110010110" => P_HR_S519 <= P_HR_S519 + T_STRESS;
				when "01110011001" => P_HR_S520 <= P_HR_S520 + T_STRESS;
				when "01110011011" => P_HR_S521 <= P_HR_S521 + T_STRESS;
				when "01110011110" => P_HR_S522 <= P_HR_S522 + T_STRESS;
				when "01110100000" => P_HR_S523 <= P_HR_S523 + T_STRESS;
				when "01110100011" => P_HR_S524 <= P_HR_S524 + T_STRESS;
				when "01110100101" => P_HR_S525 <= P_HR_S525 + T_STRESS;
				when "01110101000" => P_HR_S526 <= P_HR_S526 + T_STRESS;
				when "01110101011" => P_HR_S527 <= P_HR_S527 + T_STRESS;
				when "01110101101" => P_HR_S528 <= P_HR_S528 + T_STRESS;
				when "01110110000" => P_HR_S529 <= P_HR_S529 + T_STRESS;
				when "01110110010" => P_HR_S530 <= P_HR_S530 + T_STRESS;
				when "01110110101" => P_HR_S531 <= P_HR_S531 + T_STRESS;
				when "01110111000" => P_HR_S532 <= P_HR_S532 + T_STRESS;
				when "01110111011" => P_HR_S533 <= P_HR_S533 + T_STRESS;
				when "01110111101" => P_HR_S534 <= P_HR_S534 + T_STRESS;
				when "01111000000" => P_HR_S535 <= P_HR_S535 + T_STRESS;
				when "01111000011" => P_HR_S536 <= P_HR_S536 + T_STRESS;
				when "01111000110" => P_HR_S537 <= P_HR_S537 + T_STRESS;
				when "01111001000" => P_HR_S538 <= P_HR_S538 + T_STRESS;
				when "01111001011" => P_HR_S539 <= P_HR_S539 + T_STRESS;
				when "01111001110" => P_HR_S540 <= P_HR_S540 + T_STRESS;
				when "01111010001" => P_HR_S541 <= P_HR_S541 + T_STRESS;
				when "01111010100" => P_HR_S542 <= P_HR_S542 + T_STRESS;
				when "01111010110" => P_HR_S543 <= P_HR_S543 + T_STRESS;
				when "01111011001" => P_HR_S544 <= P_HR_S544 + T_STRESS;
				when "01111011100" => P_HR_S545 <= P_HR_S545 + T_STRESS;
				when "01111011111" => P_HR_S546 <= P_HR_S546 + T_STRESS;
				when "01111100010" => P_HR_S547 <= P_HR_S547 + T_STRESS;
				when "01111100101" => P_HR_S548 <= P_HR_S548 + T_STRESS;
				when "01111101000" => P_HR_S549 <= P_HR_S549 + T_STRESS;
				when "01111101011" => P_HR_S550 <= P_HR_S550 + T_STRESS;
				when "01111101110" => P_HR_S551 <= P_HR_S551 + T_STRESS;
				when "01111110001" => P_HR_S552 <= P_HR_S552 + T_STRESS;
				when "01111110100" => P_HR_S553 <= P_HR_S553 + T_STRESS;
				when "01111110111" => P_HR_S554 <= P_HR_S554 + T_STRESS;
				when "01111111010" => P_HR_S555 <= P_HR_S555 + T_STRESS;
				when "01111111101" => P_HR_S556 <= P_HR_S556 + T_STRESS;
				when "10000000000" => P_HR_S557 <= P_HR_S557 + T_STRESS;
				when "10000000100" => P_HR_S558 <= P_HR_S558 + T_STRESS;
				when "10000000111" => P_HR_S559 <= P_HR_S559 + T_STRESS;
				when "10000001010" => P_HR_S560 <= P_HR_S560 + T_STRESS;
				when "10000001101" => P_HR_S561 <= P_HR_S561 + T_STRESS;
				when "10000010000" => P_HR_S562 <= P_HR_S562 + T_STRESS;
				when "10000010011" => P_HR_S563 <= P_HR_S563 + T_STRESS;
				when "10000010111" => P_HR_S564 <= P_HR_S564 + T_STRESS;
				when "10000011010" => P_HR_S565 <= P_HR_S565 + T_STRESS;
				when "10000011101" => P_HR_S566 <= P_HR_S566 + T_STRESS;
				when "10000100001" => P_HR_S567 <= P_HR_S567 + T_STRESS;
				when "10000100100" => P_HR_S568 <= P_HR_S568 + T_STRESS;
				when "10000100111" => P_HR_S569 <= P_HR_S569 + T_STRESS;
				when "10000101011" => P_HR_S570 <= P_HR_S570 + T_STRESS;
				when "10000101110" => P_HR_S571 <= P_HR_S571 + T_STRESS;
				when "10000110001" => P_HR_S572 <= P_HR_S572 + T_STRESS;
				when "10000110101" => P_HR_S573 <= P_HR_S573 + T_STRESS;
				when "10000111000" => P_HR_S574 <= P_HR_S574 + T_STRESS;
				when "10000111100" => P_HR_S575 <= P_HR_S575 + T_STRESS;
				when "10000111111" => P_HR_S576 <= P_HR_S576 + T_STRESS;
				when "10001000011" => P_HR_S577 <= P_HR_S577 + T_STRESS;
				when "10001000110" => P_HR_S578 <= P_HR_S578 + T_STRESS;
				when "10001001010" => P_HR_S579 <= P_HR_S579 + T_STRESS;
				when "10001001110" => P_HR_S580 <= P_HR_S580 + T_STRESS;
				when "10001010001" => P_HR_S581 <= P_HR_S581 + T_STRESS;
				when "10001010101" => P_HR_S582 <= P_HR_S582 + T_STRESS;
				when "10001011001" => P_HR_S583 <= P_HR_S583 + T_STRESS;
				when "10001011100" => P_HR_S584 <= P_HR_S584 + T_STRESS;
				when "10001100000" => P_HR_S585 <= P_HR_S585 + T_STRESS;
				when "10001100100" => P_HR_S586 <= P_HR_S586 + T_STRESS;
				when "10001101000" => P_HR_S587 <= P_HR_S587 + T_STRESS;
				when "10001101011" => P_HR_S588 <= P_HR_S588 + T_STRESS;
				when "10001101111" => P_HR_S589 <= P_HR_S589 + T_STRESS;
				when "10001110011" => P_HR_S590 <= P_HR_S590 + T_STRESS;
				when "10001110111" => P_HR_S591 <= P_HR_S591 + T_STRESS;
				when "10001111011" => P_HR_S592 <= P_HR_S592 + T_STRESS;
				when "10001111111" => P_HR_S593 <= P_HR_S593 + T_STRESS;
				when "10010000011" => P_HR_S594 <= P_HR_S594 + T_STRESS;
				when "10010000111" => P_HR_S595 <= P_HR_S595 + T_STRESS;
				when "10010001011" => P_HR_S596 <= P_HR_S596 + T_STRESS;
				when "10010001111" => P_HR_S597 <= P_HR_S597 + T_STRESS;
				when "10010010011" => P_HR_S598 <= P_HR_S598 + T_STRESS;
				when "10010010111" => P_HR_S599 <= P_HR_S599 + T_STRESS;
				when "10010011011" => P_HR_S600 <= P_HR_S600 + T_STRESS;
				when "10010011111" => P_HR_S601 <= P_HR_S601 + T_STRESS;
				when "10010100011" => P_HR_S602 <= P_HR_S602 + T_STRESS;
				when "10010100111" => P_HR_S603 <= P_HR_S603 + T_STRESS;
				when "10010101100" => P_HR_S604 <= P_HR_S604 + T_STRESS;
				when "10010110000" => P_HR_S605 <= P_HR_S605 + T_STRESS;
				when "10010110100" => P_HR_S606 <= P_HR_S606 + T_STRESS;
				when "10010111001" => P_HR_S607 <= P_HR_S607 + T_STRESS;
				when "10010111101" => P_HR_S608 <= P_HR_S608 + T_STRESS;
				when "10011000001" => P_HR_S609 <= P_HR_S609 + T_STRESS;
				when "10011000110" => P_HR_S610 <= P_HR_S610 + T_STRESS;
				when "10011001010" => P_HR_S611 <= P_HR_S611 + T_STRESS;
				when "10011001111" => P_HR_S612 <= P_HR_S612 + T_STRESS;
				when "10011010011" => P_HR_S613 <= P_HR_S613 + T_STRESS;
				when "10011011000" => P_HR_S614 <= P_HR_S614 + T_STRESS;
				when "10011011100" => P_HR_S615 <= P_HR_S615 + T_STRESS;
				when "10011100001" => P_HR_S616 <= P_HR_S616 + T_STRESS;
				when "10011100110" => P_HR_S617 <= P_HR_S617 + T_STRESS;
				when "10011101010" => P_HR_S618 <= P_HR_S618 + T_STRESS;
				when "10011101111" => P_HR_S619 <= P_HR_S619 + T_STRESS;
				when "10100000010" => P_HR_S620 <= P_HR_S620 + T_STRESS;
				when "10100100110" => P_HR_S621 <= P_HR_S621 + T_STRESS;
				when "11001101111" => P_HR_S622 <= P_HR_S622 + T_STRESS;
				when "11010110010" => P_HR_S623 <= P_HR_S623 + T_STRESS;
				when "11011011111" => P_HR_S624 <= P_HR_S624 + T_STRESS;
				when others            => null;
			end case;

			case eda is
				when "00001000" => P_EDA_S1 <= P_EDA_S1 + T_STRESS;
				when "00001001" => P_EDA_S2 <= P_EDA_S2 + T_STRESS;
				when "00001010" => P_EDA_S3 <= P_EDA_S3 + T_STRESS;
				when "00001011" => P_EDA_S4 <= P_EDA_S4 + T_STRESS;
				when "00001100" => P_EDA_S5 <= P_EDA_S5 + T_STRESS;
				when "00001101" => P_EDA_S6 <= P_EDA_S6 + T_STRESS;
				when "00001110" => P_EDA_S7 <= P_EDA_S7 + T_STRESS;
				when "00001111" => P_EDA_S8 <= P_EDA_S8 + T_STRESS;
				when "00010000" => P_EDA_S9 <= P_EDA_S9 + T_STRESS;
				when "00010001" => P_EDA_S10 <= P_EDA_S10 + T_STRESS;
				when "00010010" => P_EDA_S11 <= P_EDA_S11 + T_STRESS;
				when "00010011" => P_EDA_S12 <= P_EDA_S12 + T_STRESS;
				when "00010100" => P_EDA_S13 <= P_EDA_S13 + T_STRESS;
				when "00010101" => P_EDA_S14 <= P_EDA_S14 + T_STRESS;
				when "00010110" => P_EDA_S15 <= P_EDA_S15 + T_STRESS;
				when "00010111" => P_EDA_S16 <= P_EDA_S16 + T_STRESS;
				when "00011000" => P_EDA_S17 <= P_EDA_S17 + T_STRESS;
				when "00011001" => P_EDA_S18 <= P_EDA_S18 + T_STRESS;
				when "00011010" => P_EDA_S19 <= P_EDA_S19 + T_STRESS;
				when "00011011" => P_EDA_S20 <= P_EDA_S20 + T_STRESS;
				when "00011100" => P_EDA_S21 <= P_EDA_S21 + T_STRESS;
				when "00011101" => P_EDA_S22 <= P_EDA_S22 + T_STRESS;
				when "00011110" => P_EDA_S23 <= P_EDA_S23 + T_STRESS;
				when "00011111" => P_EDA_S24 <= P_EDA_S24 + T_STRESS;
				when "00100000" => P_EDA_S25 <= P_EDA_S25 + T_STRESS;
				when "00100001" => P_EDA_S26 <= P_EDA_S26 + T_STRESS;
				when "00100010" => P_EDA_S27 <= P_EDA_S27 + T_STRESS;
				when "00100011" => P_EDA_S28 <= P_EDA_S28 + T_STRESS;
				when "00100100" => P_EDA_S29 <= P_EDA_S29 + T_STRESS;
				when "00100101" => P_EDA_S30 <= P_EDA_S30 + T_STRESS;
				when "00100110" => P_EDA_S31 <= P_EDA_S31 + T_STRESS;
				when "00100111" => P_EDA_S32 <= P_EDA_S32 + T_STRESS;
				when "00101000" => P_EDA_S33 <= P_EDA_S33 + T_STRESS;
				when "00101001" => P_EDA_S34 <= P_EDA_S34 + T_STRESS;
				when "00101010" => P_EDA_S35 <= P_EDA_S35 + T_STRESS;
				when "00101011" => P_EDA_S36 <= P_EDA_S36 + T_STRESS;
				when "00101100" => P_EDA_S37 <= P_EDA_S37 + T_STRESS;
				when "00101101" => P_EDA_S38 <= P_EDA_S38 + T_STRESS;
				when "00101110" => P_EDA_S39 <= P_EDA_S39 + T_STRESS;
				when "00101111" => P_EDA_S40 <= P_EDA_S40 + T_STRESS;
				when "00110000" => P_EDA_S41 <= P_EDA_S41 + T_STRESS;
				when "00110001" => P_EDA_S42 <= P_EDA_S42 + T_STRESS;
				when "00110010" => P_EDA_S43 <= P_EDA_S43 + T_STRESS;
				when "00110011" => P_EDA_S44 <= P_EDA_S44 + T_STRESS;
				when "00110100" => P_EDA_S45 <= P_EDA_S45 + T_STRESS;
				when "00110101" => P_EDA_S46 <= P_EDA_S46 + T_STRESS;
				when "00110110" => P_EDA_S47 <= P_EDA_S47 + T_STRESS;
				when "00110111" => P_EDA_S48 <= P_EDA_S48 + T_STRESS;
				when "00111000" => P_EDA_S49 <= P_EDA_S49 + T_STRESS;
				when "00111001" => P_EDA_S50 <= P_EDA_S50 + T_STRESS;
				when "00111010" => P_EDA_S51 <= P_EDA_S51 + T_STRESS;
				when "00111011" => P_EDA_S52 <= P_EDA_S52 + T_STRESS;
				when "00111100" => P_EDA_S53 <= P_EDA_S53 + T_STRESS;
				when "00111101" => P_EDA_S54 <= P_EDA_S54 + T_STRESS;
				when "00111110" => P_EDA_S55 <= P_EDA_S55 + T_STRESS;
				when "00111111" => P_EDA_S56 <= P_EDA_S56 + T_STRESS;
				when "01000000" => P_EDA_S57 <= P_EDA_S57 + T_STRESS;
				when "01000001" => P_EDA_S58 <= P_EDA_S58 + T_STRESS;
				when "01000010" => P_EDA_S59 <= P_EDA_S59 + T_STRESS;
				when "01000011" => P_EDA_S60 <= P_EDA_S60 + T_STRESS;
				when "01000100" => P_EDA_S61 <= P_EDA_S61 + T_STRESS;
				when "01000101" => P_EDA_S62 <= P_EDA_S62 + T_STRESS;
				when "01000110" => P_EDA_S63 <= P_EDA_S63 + T_STRESS;
				when "01000111" => P_EDA_S64 <= P_EDA_S64 + T_STRESS;
				when "01001000" => P_EDA_S65 <= P_EDA_S65 + T_STRESS;
				when "01001001" => P_EDA_S66 <= P_EDA_S66 + T_STRESS;
				when "01001010" => P_EDA_S67 <= P_EDA_S67 + T_STRESS;
				when "01001011" => P_EDA_S68 <= P_EDA_S68 + T_STRESS;
				when "01001100" => P_EDA_S69 <= P_EDA_S69 + T_STRESS;
				when "01001101" => P_EDA_S70 <= P_EDA_S70 + T_STRESS;
				when "01001110" => P_EDA_S71 <= P_EDA_S71 + T_STRESS;
				when "01001111" => P_EDA_S72 <= P_EDA_S72 + T_STRESS;
				when "01010000" => P_EDA_S73 <= P_EDA_S73 + T_STRESS;
				when "01010001" => P_EDA_S74 <= P_EDA_S74 + T_STRESS;
				when "01010010" => P_EDA_S75 <= P_EDA_S75 + T_STRESS;
				when "01010011" => P_EDA_S76 <= P_EDA_S76 + T_STRESS;
				when "01010100" => P_EDA_S77 <= P_EDA_S77 + T_STRESS;
				when "01010101" => P_EDA_S78 <= P_EDA_S78 + T_STRESS;
				when "01010110" => P_EDA_S79 <= P_EDA_S79 + T_STRESS;
				when "01010111" => P_EDA_S80 <= P_EDA_S80 + T_STRESS;
				when "01011000" => P_EDA_S81 <= P_EDA_S81 + T_STRESS;
				when "01011001" => P_EDA_S82 <= P_EDA_S82 + T_STRESS;
				when "01011010" => P_EDA_S83 <= P_EDA_S83 + T_STRESS;
				when "01011011" => P_EDA_S84 <= P_EDA_S84 + T_STRESS;
				when "01011100" => P_EDA_S85 <= P_EDA_S85 + T_STRESS;
				when "01011101" => P_EDA_S86 <= P_EDA_S86 + T_STRESS;
				when "01011110" => P_EDA_S87 <= P_EDA_S87 + T_STRESS;
				when "01011111" => P_EDA_S88 <= P_EDA_S88 + T_STRESS;
				when "01100000" => P_EDA_S89 <= P_EDA_S89 + T_STRESS;
				when "01100001" => P_EDA_S90 <= P_EDA_S90 + T_STRESS;
				when "01111001" => P_EDA_S91 <= P_EDA_S91 + T_STRESS;
				when "01111010" => P_EDA_S92 <= P_EDA_S92 + T_STRESS;
				when "01111011" => P_EDA_S93 <= P_EDA_S93 + T_STRESS;
				when "01111100" => P_EDA_S94 <= P_EDA_S94 + T_STRESS;
				when "01111101" => P_EDA_S95 <= P_EDA_S95 + T_STRESS;
				when "01111110" => P_EDA_S96 <= P_EDA_S96 + T_STRESS;
				when "01111111" => P_EDA_S97 <= P_EDA_S97 + T_STRESS;
				when "10000000" => P_EDA_S98 <= P_EDA_S98 + T_STRESS;
				when "10000001" => P_EDA_S99 <= P_EDA_S99 + T_STRESS;
				when "10000010" => P_EDA_S100 <= P_EDA_S100 + T_STRESS;
				when "10000011" => P_EDA_S101 <= P_EDA_S101 + T_STRESS;
				when "10000100" => P_EDA_S102 <= P_EDA_S102 + T_STRESS;
				when "10000101" => P_EDA_S103 <= P_EDA_S103 + T_STRESS;
				when "10000110" => P_EDA_S104 <= P_EDA_S104 + T_STRESS;
				when "10000111" => P_EDA_S105 <= P_EDA_S105 + T_STRESS;
				when "10001000" => P_EDA_S106 <= P_EDA_S106 + T_STRESS;
				when "10001001" => P_EDA_S107 <= P_EDA_S107 + T_STRESS;
				when "10001010" => P_EDA_S108 <= P_EDA_S108 + T_STRESS;
				when "10001011" => P_EDA_S109 <= P_EDA_S109 + T_STRESS;
				when "10001100" => P_EDA_S110 <= P_EDA_S110 + T_STRESS;
				when "10001101" => P_EDA_S111 <= P_EDA_S111 + T_STRESS;
				when "10001110" => P_EDA_S112 <= P_EDA_S112 + T_STRESS;
				when "10001111" => P_EDA_S113 <= P_EDA_S113 + T_STRESS;
				when "10010000" => P_EDA_S114 <= P_EDA_S114 + T_STRESS;
				when "10010001" => P_EDA_S115 <= P_EDA_S115 + T_STRESS;
				when "10010010" => P_EDA_S116 <= P_EDA_S116 + T_STRESS;
				when "10010011" => P_EDA_S117 <= P_EDA_S117 + T_STRESS;
				when "10010100" => P_EDA_S118 <= P_EDA_S118 + T_STRESS;
				when "10010101" => P_EDA_S119 <= P_EDA_S119 + T_STRESS;
				when "10010110" => P_EDA_S120 <= P_EDA_S120 + T_STRESS;
				when "10010111" => P_EDA_S121 <= P_EDA_S121 + T_STRESS;
				when "10011000" => P_EDA_S122 <= P_EDA_S122 + T_STRESS;
				when "10011001" => P_EDA_S123 <= P_EDA_S123 + T_STRESS;
				when "10011010" => P_EDA_S124 <= P_EDA_S124 + T_STRESS;
				when "10011011" => P_EDA_S125 <= P_EDA_S125 + T_STRESS;
				when "10011100" => P_EDA_S126 <= P_EDA_S126 + T_STRESS;
				when "10011101" => P_EDA_S127 <= P_EDA_S127 + T_STRESS;
				when "10011110" => P_EDA_S128 <= P_EDA_S128 + T_STRESS;
				when "10011111" => P_EDA_S129 <= P_EDA_S129 + T_STRESS;
				when "10100000" => P_EDA_S130 <= P_EDA_S130 + T_STRESS;
				when others            => null;
			end case;
		    
		else -- not in normal or training mode
			stress_score <= (others => '0');
			P_TEMP_S <= (others => '0'); 
			P_EDA_S <= (others => '0');
			P_HR_S <= (others => '0');
		end if;
		end if;
	end process;
	
	process(clk, rst) -- not stressed
	begin
	if (rst = '1') then
		-- reset logic
        P_TEMP_NS1 <= (others => '0');
        P_TEMP_NS2 <= (others => '0');
        P_TEMP_NS3 <= (others => '0');
        P_TEMP_NS4 <= (others => '0');
        P_TEMP_NS5 <= (others => '0');
        P_TEMP_NS6 <= (others => '0');
        P_TEMP_NS7 <= (others => '0');
        P_TEMP_NS8 <= (others => '0');
        P_TEMP_NS9 <= (others => '0');
        P_TEMP_NS10 <= (others => '0');
        P_TEMP_NS11 <= (others => '0');
        P_TEMP_NS12 <= (others => '0');
        P_TEMP_NS13 <= (others => '0');
        P_TEMP_NS14 <= (others => '0');
        P_TEMP_NS15 <= (others => '0');
        P_TEMP_NS16 <= (others => '0');
        P_TEMP_NS17 <= (others => '0');
        P_TEMP_NS18 <= (others => '0');
        P_TEMP_NS19 <= (others => '0');
        P_TEMP_NS20 <= (others => '0');
        P_TEMP_NS21 <= (others => '0');
        P_TEMP_NS22 <= (others => '0');
        P_TEMP_NS23 <= (others => '0');
        P_TEMP_NS24 <= (others => '0');
        P_TEMP_NS25 <= (others => '0');
        P_TEMP_NS26 <= (others => '0');
        P_TEMP_NS27 <= (others => '0');
        P_TEMP_NS28 <= (others => '0');
        P_TEMP_NS29 <= (others => '0');
        P_TEMP_NS30 <= (others => '0');
        P_TEMP_NS31 <= (others => '0');
        P_TEMP_NS32 <= (others => '0');
        P_TEMP_NS33 <= (others => '0');
        P_TEMP_NS34 <= (others => '0');
        P_TEMP_NS35 <= (others => '0');
        P_TEMP_NS36 <= (others => '0');
        P_TEMP_NS37 <= (others => '0');
        P_TEMP_NS38 <= (others => '0');
        P_TEMP_NS39 <= (others => '0');
        P_TEMP_NS40 <= (others => '0');
        P_TEMP_NS41 <= (others => '0');
        P_TEMP_NS42 <= (others => '0');
        P_TEMP_NS43 <= (others => '0');
        P_TEMP_NS44 <= (others => '0');
        P_TEMP_NS45 <= (others => '0');
        P_TEMP_NS46 <= (others => '0');
        P_TEMP_NS47 <= (others => '0');
        P_TEMP_NS48 <= (others => '0');
        P_TEMP_NS49 <= (others => '0');
        P_TEMP_NS50 <= (others => '0');
        P_TEMP_NS51 <= (others => '0');
        P_TEMP_NS52 <= (others => '0');
        P_TEMP_NS53 <= (others => '0');
        P_TEMP_NS54 <= (others => '0');
        P_TEMP_NS55 <= (others => '0');
        P_TEMP_NS56 <= (others => '0');
        P_TEMP_NS57 <= (others => '0');
        P_TEMP_NS58 <= (others => '0');
        P_TEMP_NS59 <= (others => '0');
        P_TEMP_NS60 <= (others => '0');
        P_TEMP_NS61 <= (others => '0');
        P_TEMP_NS62 <= (others => '0');
        P_TEMP_NS63 <= (others => '0');
			
        P_HR_NS1 <= (others => '0');
        P_HR_NS2 <= (others => '0');
        P_HR_NS3 <= (others => '0');
        P_HR_NS4 <= (others => '0');
        P_HR_NS5 <= (others => '0');
        P_HR_NS6 <= (others => '0');
        P_HR_NS7 <= (others => '0');
        P_HR_NS8 <= (others => '0');
        P_HR_NS9 <= (others => '0');
        P_HR_NS10 <= (others => '0');
        P_HR_NS11 <= (others => '0');
        P_HR_NS12 <= (others => '0');
        P_HR_NS13 <= (others => '0');
        P_HR_NS14 <= (others => '0');
        P_HR_NS15 <= (others => '0');
        P_HR_NS16 <= (others => '0');
        P_HR_NS17 <= (others => '0');
        P_HR_NS18 <= (others => '0');
        P_HR_NS19 <= (others => '0');
        P_HR_NS20 <= (others => '0');
        P_HR_NS21 <= (others => '0');
        P_HR_NS22 <= (others => '0');
        P_HR_NS23 <= (others => '0');
        P_HR_NS24 <= (others => '0');
        P_HR_NS25 <= (others => '0');
        P_HR_NS26 <= (others => '0');
        P_HR_NS27 <= (others => '0');
        P_HR_NS28 <= (others => '0');
        P_HR_NS29 <= (others => '0');
        P_HR_NS30 <= (others => '0');
        P_HR_NS31 <= (others => '0');
        P_HR_NS32 <= (others => '0');
        P_HR_NS33 <= (others => '0');
        P_HR_NS34 <= (others => '0');
        P_HR_NS35 <= (others => '0');
        P_HR_NS36 <= (others => '0');
        P_HR_NS37 <= (others => '0');
        P_HR_NS38 <= (others => '0');
        P_HR_NS39 <= (others => '0');
        P_HR_NS40 <= (others => '0');
        P_HR_NS41 <= (others => '0');
        P_HR_NS42 <= (others => '0');
        P_HR_NS43 <= (others => '0');
        P_HR_NS44 <= (others => '0');
        P_HR_NS45 <= (others => '0');
        P_HR_NS46 <= (others => '0');
        P_HR_NS47 <= (others => '0');
        P_HR_NS48 <= (others => '0');
        P_HR_NS49 <= (others => '0');
        P_HR_NS50 <= (others => '0');
        P_HR_NS51 <= (others => '0');
        P_HR_NS52 <= (others => '0');
        P_HR_NS53 <= (others => '0');
        P_HR_NS54 <= (others => '0');
        P_HR_NS55 <= (others => '0');
        P_HR_NS56 <= (others => '0');
        P_HR_NS57 <= (others => '0');
        P_HR_NS58 <= (others => '0');
        P_HR_NS59 <= (others => '0');
        P_HR_NS60 <= (others => '0');
        P_HR_NS61 <= (others => '0');
        P_HR_NS62 <= (others => '0');
        P_HR_NS63 <= (others => '0');
        P_HR_NS64 <= (others => '0');
        P_HR_NS65 <= (others => '0');
        P_HR_NS66 <= (others => '0');
        P_HR_NS67 <= (others => '0');
        P_HR_NS68 <= (others => '0');
        P_HR_NS69 <= (others => '0');
        P_HR_NS70 <= (others => '0');
        P_HR_NS71 <= (others => '0');
        P_HR_NS72 <= (others => '0');
        P_HR_NS73 <= (others => '0');
        P_HR_NS74 <= (others => '0');
        P_HR_NS75 <= (others => '0');
        P_HR_NS76 <= (others => '0');
        P_HR_NS77 <= (others => '0');
        P_HR_NS78 <= (others => '0');
        P_HR_NS79 <= (others => '0');
        P_HR_NS80 <= (others => '0');
        P_HR_NS81 <= (others => '0');
        P_HR_NS82 <= (others => '0');
        P_HR_NS83 <= (others => '0');
        P_HR_NS84 <= (others => '0');
        P_HR_NS85 <= (others => '0');
        P_HR_NS86 <= (others => '0');
        P_HR_NS87 <= (others => '0');
        P_HR_NS88 <= (others => '0');
        P_HR_NS89 <= (others => '0');
        P_HR_NS90 <= (others => '0');
        P_HR_NS91 <= (others => '0');
        P_HR_NS92 <= (others => '0');
        P_HR_NS93 <= (others => '0');
        P_HR_NS94 <= (others => '0');
        P_HR_NS95 <= (others => '0');
        P_HR_NS96 <= (others => '0');
        P_HR_NS97 <= (others => '0');
        P_HR_NS98 <= (others => '0');
        P_HR_NS99 <= (others => '0');
        P_HR_NS100 <= (others => '0');
        P_HR_NS101 <= (others => '0');
        P_HR_NS102 <= (others => '0');
        P_HR_NS103 <= (others => '0');
        P_HR_NS104 <= (others => '0');
        P_HR_NS105 <= (others => '0');
        P_HR_NS106 <= (others => '0');
        P_HR_NS107 <= (others => '0');
        P_HR_NS108 <= (others => '0');
        P_HR_NS109 <= (others => '0');
        P_HR_NS110 <= (others => '0');
        P_HR_NS111 <= (others => '0');
        P_HR_NS112 <= (others => '0');
        P_HR_NS113 <= (others => '0');
        P_HR_NS114 <= (others => '0');
        P_HR_NS115 <= (others => '0');
        P_HR_NS116 <= (others => '0');
        P_HR_NS117 <= (others => '0');
        P_HR_NS118 <= (others => '0');
        P_HR_NS119 <= (others => '0');
        P_HR_NS120 <= (others => '0');
        P_HR_NS121 <= (others => '0');
        P_HR_NS122 <= (others => '0');
        P_HR_NS123 <= (others => '0');
        P_HR_NS124 <= (others => '0');
        P_HR_NS125 <= (others => '0');
        P_HR_NS126 <= (others => '0');
        P_HR_NS127 <= (others => '0');
        P_HR_NS128 <= (others => '0');
        P_HR_NS129 <= (others => '0');
        P_HR_NS130 <= (others => '0');
        P_HR_NS131 <= (others => '0');
        P_HR_NS132 <= (others => '0');
        P_HR_NS133 <= (others => '0');
        P_HR_NS134 <= (others => '0');
        P_HR_NS135 <= (others => '0');
        P_HR_NS136 <= (others => '0');
        P_HR_NS137 <= (others => '0');
        P_HR_NS138 <= (others => '0');
        P_HR_NS139 <= (others => '0');
        P_HR_NS140 <= (others => '0');
        P_HR_NS141 <= (others => '0');
        P_HR_NS142 <= (others => '0');
        P_HR_NS143 <= (others => '0');
        P_HR_NS144 <= (others => '0');
        P_HR_NS145 <= (others => '0');
        P_HR_NS146 <= (others => '0');
        P_HR_NS147 <= (others => '0');
        P_HR_NS148 <= (others => '0');
        P_HR_NS149 <= (others => '0');
        P_HR_NS150 <= (others => '0');
        P_HR_NS151 <= (others => '0');
        P_HR_NS152 <= (others => '0');
        P_HR_NS153 <= (others => '0');
        P_HR_NS154 <= (others => '0');
        P_HR_NS155 <= (others => '0');
        P_HR_NS156 <= (others => '0');
        P_HR_NS157 <= (others => '0');
        P_HR_NS158 <= (others => '0');
        P_HR_NS159 <= (others => '0');
        P_HR_NS160 <= (others => '0');
        P_HR_NS161 <= (others => '0');
        P_HR_NS162 <= (others => '0');
        P_HR_NS163 <= (others => '0');
        P_HR_NS164 <= (others => '0');
        P_HR_NS165 <= (others => '0');
        P_HR_NS166 <= (others => '0');
        P_HR_NS167 <= (others => '0');
        P_HR_NS168 <= (others => '0');
        P_HR_NS169 <= (others => '0');
        P_HR_NS170 <= (others => '0');
        P_HR_NS171 <= (others => '0');
        P_HR_NS172 <= (others => '0');
        P_HR_NS173 <= (others => '0');
        P_HR_NS174 <= (others => '0');
        P_HR_NS175 <= (others => '0');
        P_HR_NS176 <= (others => '0');
        P_HR_NS177 <= (others => '0');
        P_HR_NS178 <= (others => '0');
        P_HR_NS179 <= (others => '0');
        P_HR_NS180 <= (others => '0');
        P_HR_NS181 <= (others => '0');
        P_HR_NS182 <= (others => '0');
        P_HR_NS183 <= (others => '0');
        P_HR_NS184 <= (others => '0');
        P_HR_NS185 <= (others => '0');
        P_HR_NS186 <= (others => '0');
        P_HR_NS187 <= (others => '0');
        P_HR_NS188 <= (others => '0');
        P_HR_NS189 <= (others => '0');
        P_HR_NS190 <= (others => '0');
        P_HR_NS191 <= (others => '0');
        P_HR_NS192 <= (others => '0');
        P_HR_NS193 <= (others => '0');
        P_HR_NS194 <= (others => '0');
        P_HR_NS195 <= (others => '0');
        P_HR_NS196 <= (others => '0');
        P_HR_NS197 <= (others => '0');
        P_HR_NS198 <= (others => '0');
        P_HR_NS199 <= (others => '0');
        P_HR_NS200 <= (others => '0');
        P_HR_NS201 <= (others => '0');
        P_HR_NS202 <= (others => '0');
        P_HR_NS203 <= (others => '0');
        P_HR_NS204 <= (others => '0');
        P_HR_NS205 <= (others => '0');
        P_HR_NS206 <= (others => '0');
        P_HR_NS207 <= (others => '0');
        P_HR_NS208 <= (others => '0');
        P_HR_NS209 <= (others => '0');
        P_HR_NS210 <= (others => '0');
        P_HR_NS211 <= (others => '0');
        P_HR_NS212 <= (others => '0');
        P_HR_NS213 <= (others => '0');
        P_HR_NS214 <= (others => '0');
        P_HR_NS215 <= (others => '0');
        P_HR_NS216 <= (others => '0');
        P_HR_NS217 <= (others => '0');
        P_HR_NS218 <= (others => '0');
        P_HR_NS219 <= (others => '0');
        P_HR_NS220 <= (others => '0');
        P_HR_NS221 <= (others => '0');
        P_HR_NS222 <= (others => '0');
        P_HR_NS223 <= (others => '0');
        P_HR_NS224 <= (others => '0');
        P_HR_NS225 <= (others => '0');
        P_HR_NS226 <= (others => '0');
        P_HR_NS227 <= (others => '0');
        P_HR_NS228 <= (others => '0');
        P_HR_NS229 <= (others => '0');
        P_HR_NS230 <= (others => '0');
        P_HR_NS231 <= (others => '0');
        P_HR_NS232 <= (others => '0');
        P_HR_NS233 <= (others => '0');
        P_HR_NS234 <= (others => '0');
        P_HR_NS235 <= (others => '0');
        P_HR_NS236 <= (others => '0');
        P_HR_NS237 <= (others => '0');
        P_HR_NS238 <= (others => '0');
        P_HR_NS239 <= (others => '0');
        P_HR_NS240 <= (others => '0');
        P_HR_NS241 <= (others => '0');
        P_HR_NS242 <= (others => '0');
        P_HR_NS243 <= (others => '0');
        P_HR_NS244 <= (others => '0');
        P_HR_NS245 <= (others => '0');
        P_HR_NS246 <= (others => '0');
        P_HR_NS247 <= (others => '0');
        P_HR_NS248 <= (others => '0');
        P_HR_NS249 <= (others => '0');
        P_HR_NS250 <= (others => '0');
        P_HR_NS251 <= (others => '0');
        P_HR_NS252 <= (others => '0');
        P_HR_NS253 <= (others => '0');
        P_HR_NS254 <= (others => '0');
        P_HR_NS255 <= (others => '0');
        P_HR_NS256 <= (others => '0');
        P_HR_NS257 <= (others => '0');
        P_HR_NS258 <= (others => '0');
        P_HR_NS259 <= (others => '0');
        P_HR_NS260 <= (others => '0');
        P_HR_NS261 <= (others => '0');
        P_HR_NS262 <= (others => '0');
        P_HR_NS263 <= (others => '0');
        P_HR_NS264 <= (others => '0');
        P_HR_NS265 <= (others => '0');
        P_HR_NS266 <= (others => '0');
        P_HR_NS267 <= (others => '0');
        P_HR_NS268 <= (others => '0');
        P_HR_NS269 <= (others => '0');
        P_HR_NS270 <= (others => '0');
        P_HR_NS271 <= (others => '0');
        P_HR_NS272 <= (others => '0');
        P_HR_NS273 <= (others => '0');
        P_HR_NS274 <= (others => '0');
        P_HR_NS275 <= (others => '0');
        P_HR_NS276 <= (others => '0');
        P_HR_NS277 <= (others => '0');
        P_HR_NS278 <= (others => '0');
        P_HR_NS279 <= (others => '0');
        P_HR_NS280 <= (others => '0');
        P_HR_NS281 <= (others => '0');
        P_HR_NS282 <= (others => '0');
        P_HR_NS283 <= (others => '0');
        P_HR_NS284 <= (others => '0');
        P_HR_NS285 <= (others => '0');
        P_HR_NS286 <= (others => '0');
        P_HR_NS287 <= (others => '0');
        P_HR_NS288 <= (others => '0');
        P_HR_NS289 <= (others => '0');
        P_HR_NS290 <= (others => '0');
        P_HR_NS291 <= (others => '0');
        P_HR_NS292 <= (others => '0');
        P_HR_NS293 <= (others => '0');
        P_HR_NS294 <= (others => '0');
        P_HR_NS295 <= (others => '0');
        P_HR_NS296 <= (others => '0');
        P_HR_NS297 <= (others => '0');
        P_HR_NS298 <= (others => '0');
        P_HR_NS299 <= (others => '0');
        P_HR_NS300 <= (others => '0');
        P_HR_NS301 <= (others => '0');
        P_HR_NS302 <= (others => '0');
        P_HR_NS303 <= (others => '0');
        P_HR_NS304 <= (others => '0');
        P_HR_NS305 <= (others => '0');
        P_HR_NS306 <= (others => '0');
        P_HR_NS307 <= (others => '0');
        P_HR_NS308 <= (others => '0');
        P_HR_NS309 <= (others => '0');
        P_HR_NS310 <= (others => '0');
        P_HR_NS311 <= (others => '0');
        P_HR_NS312 <= (others => '0');
        P_HR_NS313 <= (others => '0');
        P_HR_NS314 <= (others => '0');
        P_HR_NS315 <= (others => '0');
        P_HR_NS316 <= (others => '0');
        P_HR_NS317 <= (others => '0');
        P_HR_NS318 <= (others => '0');
        P_HR_NS319 <= (others => '0');
        P_HR_NS320 <= (others => '0');
        P_HR_NS321 <= (others => '0');
        P_HR_NS322 <= (others => '0');
        P_HR_NS323 <= (others => '0');
        P_HR_NS324 <= (others => '0');
        P_HR_NS325 <= (others => '0');
        P_HR_NS326 <= (others => '0');
        P_HR_NS327 <= (others => '0');
        P_HR_NS328 <= (others => '0');
        P_HR_NS329 <= (others => '0');
        P_HR_NS330 <= (others => '0');
        P_HR_NS331 <= (others => '0');
        P_HR_NS332 <= (others => '0');
        P_HR_NS333 <= (others => '0');
        P_HR_NS334 <= (others => '0');
        P_HR_NS335 <= (others => '0');
        P_HR_NS336 <= (others => '0');
        P_HR_NS337 <= (others => '0');
        P_HR_NS338 <= (others => '0');
        P_HR_NS339 <= (others => '0');
        P_HR_NS340 <= (others => '0');
        P_HR_NS341 <= (others => '0');
        P_HR_NS342 <= (others => '0');
        P_HR_NS343 <= (others => '0');
        P_HR_NS344 <= (others => '0');
        P_HR_NS345 <= (others => '0');
        P_HR_NS346 <= (others => '0');
        P_HR_NS347 <= (others => '0');
        P_HR_NS348 <= (others => '0');
        P_HR_NS349 <= (others => '0');
        P_HR_NS350 <= (others => '0');
        P_HR_NS351 <= (others => '0');
        P_HR_NS352 <= (others => '0');
        P_HR_NS353 <= (others => '0');
        P_HR_NS354 <= (others => '0');
        P_HR_NS355 <= (others => '0');
        P_HR_NS356 <= (others => '0');
        P_HR_NS357 <= (others => '0');
        P_HR_NS358 <= (others => '0');
        P_HR_NS359 <= (others => '0');
        P_HR_NS360 <= (others => '0');
        P_HR_NS361 <= (others => '0');
        P_HR_NS362 <= (others => '0');
        P_HR_NS363 <= (others => '0');
        P_HR_NS364 <= (others => '0');
        P_HR_NS365 <= (others => '0');
        P_HR_NS366 <= (others => '0');
        P_HR_NS367 <= (others => '0');
        P_HR_NS368 <= (others => '0');
        P_HR_NS369 <= (others => '0');
        P_HR_NS370 <= (others => '0');
        P_HR_NS371 <= (others => '0');
        P_HR_NS372 <= (others => '0');
        P_HR_NS373 <= (others => '0');
        P_HR_NS374 <= (others => '0');
        P_HR_NS375 <= (others => '0');
        P_HR_NS376 <= (others => '0');
        P_HR_NS377 <= (others => '0');
        P_HR_NS378 <= (others => '0');
        P_HR_NS379 <= (others => '0');
        P_HR_NS380 <= (others => '0');
        P_HR_NS381 <= (others => '0');
        P_HR_NS382 <= (others => '0');
        P_HR_NS383 <= (others => '0');
        P_HR_NS384 <= (others => '0');
        P_HR_NS385 <= (others => '0');
        P_HR_NS386 <= (others => '0');
        P_HR_NS387 <= (others => '0');
        P_HR_NS388 <= (others => '0');
        P_HR_NS389 <= (others => '0');
        P_HR_NS390 <= (others => '0');
        P_HR_NS391 <= (others => '0');
        P_HR_NS392 <= (others => '0');
        P_HR_NS393 <= (others => '0');
        P_HR_NS394 <= (others => '0');
        P_HR_NS395 <= (others => '0');
        P_HR_NS396 <= (others => '0');
        P_HR_NS397 <= (others => '0');
        P_HR_NS398 <= (others => '0');
        P_HR_NS399 <= (others => '0');
        P_HR_NS400 <= (others => '0');
        P_HR_NS401 <= (others => '0');
        P_HR_NS402 <= (others => '0');
        P_HR_NS403 <= (others => '0');
        P_HR_NS404 <= (others => '0');
        P_HR_NS405 <= (others => '0');
        P_HR_NS406 <= (others => '0');
        P_HR_NS407 <= (others => '0');
        P_HR_NS408 <= (others => '0');
        P_HR_NS409 <= (others => '0');
        P_HR_NS410 <= (others => '0');
        P_HR_NS411 <= (others => '0');
        P_HR_NS412 <= (others => '0');
        P_HR_NS413 <= (others => '0');
        P_HR_NS414 <= (others => '0');
        P_HR_NS415 <= (others => '0');
        P_HR_NS416 <= (others => '0');
        P_HR_NS417 <= (others => '0');
        P_HR_NS418 <= (others => '0');
        P_HR_NS419 <= (others => '0');
        P_HR_NS420 <= (others => '0');
        P_HR_NS421 <= (others => '0');
        P_HR_NS422 <= (others => '0');
        P_HR_NS423 <= (others => '0');
        P_HR_NS424 <= (others => '0');
        P_HR_NS425 <= (others => '0');
        P_HR_NS426 <= (others => '0');
        P_HR_NS427 <= (others => '0');
        P_HR_NS428 <= (others => '0');
        P_HR_NS429 <= (others => '0');
        P_HR_NS430 <= (others => '0');
        P_HR_NS431 <= (others => '0');
        P_HR_NS432 <= (others => '0');
        P_HR_NS433 <= (others => '0');
        P_HR_NS434 <= (others => '0');
        P_HR_NS435 <= (others => '0');
        P_HR_NS436 <= (others => '0');
        P_HR_NS437 <= (others => '0');
        P_HR_NS438 <= (others => '0');
        P_HR_NS439 <= (others => '0');
        P_HR_NS440 <= (others => '0');
        P_HR_NS441 <= (others => '0');
        P_HR_NS442 <= (others => '0');
        P_HR_NS443 <= (others => '0');
        P_HR_NS444 <= (others => '0');
        P_HR_NS445 <= (others => '0');
        P_HR_NS446 <= (others => '0');
        P_HR_NS447 <= (others => '0');
        P_HR_NS448 <= (others => '0');
        P_HR_NS449 <= (others => '0');
        P_HR_NS450 <= (others => '0');
        P_HR_NS451 <= (others => '0');
        P_HR_NS452 <= (others => '0');
        P_HR_NS453 <= (others => '0');
        P_HR_NS454 <= (others => '0');
        P_HR_NS455 <= (others => '0');
        P_HR_NS456 <= (others => '0');
        P_HR_NS457 <= (others => '0');
        P_HR_NS458 <= (others => '0');
        P_HR_NS459 <= (others => '0');
        P_HR_NS460 <= (others => '0');
        P_HR_NS461 <= (others => '0');
        P_HR_NS462 <= (others => '0');
        P_HR_NS463 <= (others => '0');
        P_HR_NS464 <= (others => '0');
        P_HR_NS465 <= (others => '0');
        P_HR_NS466 <= (others => '0');
        P_HR_NS467 <= (others => '0');
        P_HR_NS468 <= (others => '0');
        P_HR_NS469 <= (others => '0');
        P_HR_NS470 <= (others => '0');
        P_HR_NS471 <= (others => '0');
        P_HR_NS472 <= (others => '0');
        P_HR_NS473 <= (others => '0');
        P_HR_NS474 <= (others => '0');
        P_HR_NS475 <= (others => '0');
        P_HR_NS476 <= (others => '0');
        P_HR_NS477 <= (others => '0');
        P_HR_NS478 <= (others => '0');
        P_HR_NS479 <= (others => '0');
        P_HR_NS480 <= (others => '0');
        P_HR_NS481 <= (others => '0');
        P_HR_NS482 <= (others => '0');
        P_HR_NS483 <= (others => '0');
        P_HR_NS484 <= (others => '0');
        P_HR_NS485 <= (others => '0');
        P_HR_NS486 <= (others => '0');
        P_HR_NS487 <= (others => '0');
        P_HR_NS488 <= (others => '0');
        P_HR_NS489 <= (others => '0');
        P_HR_NS490 <= (others => '0');
        P_HR_NS491 <= (others => '0');
        P_HR_NS492 <= (others => '0');
        P_HR_NS493 <= (others => '0');
        P_HR_NS494 <= (others => '0');
        P_HR_NS495 <= (others => '0');
        P_HR_NS496 <= (others => '0');
        P_HR_NS497 <= (others => '0');
        P_HR_NS498 <= (others => '0');
        P_HR_NS499 <= (others => '0');
        P_HR_NS500 <= (others => '0');
        P_HR_NS501 <= (others => '0');
        P_HR_NS502 <= (others => '0');
        P_HR_NS503 <= (others => '0');
        P_HR_NS504 <= (others => '0');
        P_HR_NS505 <= (others => '0');
        P_HR_NS506 <= (others => '0');
        P_HR_NS507 <= (others => '0');
        P_HR_NS508 <= (others => '0');
        P_HR_NS509 <= (others => '0');
        P_HR_NS510 <= (others => '0');
        P_HR_NS511 <= (others => '0');
        P_HR_NS512 <= (others => '0');
        P_HR_NS513 <= (others => '0');
        P_HR_NS514 <= (others => '0');
        P_HR_NS515 <= (others => '0');
        P_HR_NS516 <= (others => '0');
        P_HR_NS517 <= (others => '0');
        P_HR_NS518 <= (others => '0');
        P_HR_NS519 <= (others => '0');
        P_HR_NS520 <= (others => '0');
        P_HR_NS521 <= (others => '0');
        P_HR_NS522 <= (others => '0');
        P_HR_NS523 <= (others => '0');
        P_HR_NS524 <= (others => '0');
        P_HR_NS525 <= (others => '0');
        P_HR_NS526 <= (others => '0');
        P_HR_NS527 <= (others => '0');
        P_HR_NS528 <= (others => '0');
        P_HR_NS529 <= (others => '0');
        P_HR_NS530 <= (others => '0');
        P_HR_NS531 <= (others => '0');
        P_HR_NS532 <= (others => '0');
        P_HR_NS533 <= (others => '0');
        P_HR_NS534 <= (others => '0');
        P_HR_NS535 <= (others => '0');
        P_HR_NS536 <= (others => '0');
        P_HR_NS537 <= (others => '0');
        P_HR_NS538 <= (others => '0');
        P_HR_NS539 <= (others => '0');
        P_HR_NS540 <= (others => '0');
        P_HR_NS541 <= (others => '0');
        P_HR_NS542 <= (others => '0');
        P_HR_NS543 <= (others => '0');
        P_HR_NS544 <= (others => '0');
        P_HR_NS545 <= (others => '0');
        P_HR_NS546 <= (others => '0');
        P_HR_NS547 <= (others => '0');
        P_HR_NS548 <= (others => '0');
        P_HR_NS549 <= (others => '0');
        P_HR_NS550 <= (others => '0');
        P_HR_NS551 <= (others => '0');
        P_HR_NS552 <= (others => '0');
        P_HR_NS553 <= (others => '0');
        P_HR_NS554 <= (others => '0');
        P_HR_NS555 <= (others => '0');
        P_HR_NS556 <= (others => '0');
        P_HR_NS557 <= (others => '0');
        P_HR_NS558 <= (others => '0');
        P_HR_NS559 <= (others => '0');
        P_HR_NS560 <= (others => '0');
        P_HR_NS561 <= (others => '0');
        P_HR_NS562 <= (others => '0');
        P_HR_NS563 <= (others => '0');
        P_HR_NS564 <= (others => '0');
        P_HR_NS565 <= (others => '0');
        P_HR_NS566 <= (others => '0');
        P_HR_NS567 <= (others => '0');
        P_HR_NS568 <= (others => '0');
        P_HR_NS569 <= (others => '0');
        P_HR_NS570 <= (others => '0');
        P_HR_NS571 <= (others => '0');
        P_HR_NS572 <= (others => '0');
        P_HR_NS573 <= (others => '0');
        P_HR_NS574 <= (others => '0');
        P_HR_NS575 <= (others => '0');
        P_HR_NS576 <= (others => '0');
        P_HR_NS577 <= (others => '0');
        P_HR_NS578 <= (others => '0');
        P_HR_NS579 <= (others => '0');
        P_HR_NS580 <= (others => '0');
        P_HR_NS581 <= (others => '0');
        P_HR_NS582 <= (others => '0');
        P_HR_NS583 <= (others => '0');
        P_HR_NS584 <= (others => '0');
        P_HR_NS585 <= (others => '0');
        P_HR_NS586 <= (others => '0');
        P_HR_NS587 <= (others => '0');
        P_HR_NS588 <= (others => '0');
        P_HR_NS589 <= (others => '0');
        P_HR_NS590 <= (others => '0');
        P_HR_NS591 <= (others => '0');
        P_HR_NS592 <= (others => '0');
        P_HR_NS593 <= (others => '0');
        P_HR_NS594 <= (others => '0');
        P_HR_NS595 <= (others => '0');
        P_HR_NS596 <= (others => '0');
        P_HR_NS597 <= (others => '0');
        P_HR_NS598 <= (others => '0');
        P_HR_NS599 <= (others => '0');
        P_HR_NS600 <= (others => '0');
        P_HR_NS601 <= (others => '0');
        P_HR_NS602 <= (others => '0');
        P_HR_NS603 <= (others => '0');
        P_HR_NS604 <= (others => '0');
        P_HR_NS605 <= (others => '0');
        P_HR_NS606 <= (others => '0');
        P_HR_NS607 <= (others => '0');
        P_HR_NS608 <= (others => '0');
        P_HR_NS609 <= (others => '0');
        P_HR_NS610 <= (others => '0');
        P_HR_NS611 <= (others => '0');
        P_HR_NS612 <= (others => '0');
        P_HR_NS613 <= (others => '0');
        P_HR_NS614 <= (others => '0');
        P_HR_NS615 <= (others => '0');
        P_HR_NS616 <= (others => '0');
        P_HR_NS617 <= (others => '0');
        P_HR_NS618 <= (others => '0');
        P_HR_NS619 <= (others => '0');
        P_HR_NS620 <= (others => '0');
        P_HR_NS621 <= (others => '0');
        P_HR_NS622 <= (others => '0');
        P_HR_NS623 <= (others => '0');
        P_HR_NS624 <= (others => '0');
        P_HR_NS625 <= (others => '0');
        P_HR_NS626 <= (others => '0');
        P_HR_NS627 <= (others => '0');
        P_HR_NS628 <= (others => '0');
        P_HR_NS629 <= (others => '0');
        P_HR_NS630 <= (others => '0');
        P_HR_NS631 <= (others => '0');
        P_HR_NS632 <= (others => '0');
        P_HR_NS633 <= (others => '0');
        P_HR_NS634 <= (others => '0');
        P_HR_NS635 <= (others => '0');
        P_HR_NS636 <= (others => '0');
        P_HR_NS637 <= (others => '0');
        P_HR_NS638 <= (others => '0');
        P_HR_NS639 <= (others => '0');
        P_HR_NS640 <= (others => '0');
        P_HR_NS641 <= (others => '0');
        P_HR_NS642 <= (others => '0');
        P_HR_NS643 <= (others => '0');
        P_HR_NS644 <= (others => '0');
        P_HR_NS645 <= (others => '0');
        P_HR_NS646 <= (others => '0');
        P_HR_NS647 <= (others => '0');
        P_HR_NS648 <= (others => '0');
        P_HR_NS649 <= (others => '0');
        P_HR_NS650 <= (others => '0');
        P_HR_NS651 <= (others => '0');
        P_HR_NS652 <= (others => '0');
        P_HR_NS653 <= (others => '0');
        P_HR_NS654 <= (others => '0');
        P_HR_NS655 <= (others => '0');
        P_HR_NS656 <= (others => '0');
        P_HR_NS657 <= (others => '0');
        P_HR_NS658 <= (others => '0');
        P_HR_NS659 <= (others => '0');
        P_HR_NS660 <= (others => '0');
        P_HR_NS661 <= (others => '0');
        P_HR_NS662 <= (others => '0');
        P_HR_NS663 <= (others => '0');
        P_HR_NS664 <= (others => '0');
        P_HR_NS665 <= (others => '0');
        P_HR_NS666 <= (others => '0');
        P_HR_NS667 <= (others => '0');
        P_HR_NS668 <= (others => '0');
        P_HR_NS669 <= (others => '0');
        P_HR_NS670 <= (others => '0');
        P_HR_NS671 <= (others => '0');
        P_HR_NS672 <= (others => '0');
        P_HR_NS673 <= (others => '0');
        P_HR_NS674 <= (others => '0');
        P_HR_NS675 <= (others => '0');
        P_HR_NS676 <= (others => '0');
        P_HR_NS677 <= (others => '0');
        P_HR_NS678 <= (others => '0');
        P_HR_NS679 <= (others => '0');
        P_HR_NS680 <= (others => '0');
        P_HR_NS681 <= (others => '0');
        P_HR_NS682 <= (others => '0');
        P_HR_NS683 <= (others => '0');
        P_HR_NS684 <= (others => '0');
        P_HR_NS685 <= (others => '0');
        P_HR_NS686 <= (others => '0');
        P_HR_NS687 <= (others => '0');
        P_HR_NS688 <= (others => '0');
        P_HR_NS689 <= (others => '0');
        P_HR_NS690 <= (others => '0');
        P_HR_NS691 <= (others => '0');
        P_HR_NS692 <= (others => '0');
        P_HR_NS693 <= (others => '0');
        P_HR_NS694 <= (others => '0');
        P_HR_NS695 <= (others => '0');
        P_HR_NS696 <= (others => '0');
        P_HR_NS697 <= (others => '0');
        P_HR_NS698 <= (others => '0');
        P_HR_NS699 <= (others => '0');
        P_HR_NS700 <= (others => '0');
        P_HR_NS701 <= (others => '0');
        P_HR_NS702 <= (others => '0');
        P_HR_NS703 <= (others => '0');
        P_HR_NS704 <= (others => '0');
        P_HR_NS705 <= (others => '0');
        P_HR_NS706 <= (others => '0');
        P_HR_NS707 <= (others => '0');
        P_HR_NS708 <= (others => '0');
        P_HR_NS709 <= (others => '0');
        P_HR_NS710 <= (others => '0');
        P_HR_NS711 <= (others => '0');
        P_HR_NS712 <= (others => '0');
        P_HR_NS713 <= (others => '0');
        P_HR_NS714 <= (others => '0');
        P_HR_NS715 <= (others => '0');
        P_HR_NS716 <= (others => '0');
        P_HR_NS717 <= (others => '0');
        P_HR_NS718 <= (others => '0');
        P_HR_NS719 <= (others => '0');
        P_HR_NS720 <= (others => '0');
        P_HR_NS721 <= (others => '0');
        P_HR_NS722 <= (others => '0');
        P_HR_NS723 <= (others => '0');
        P_HR_NS724 <= (others => '0');
        P_HR_NS725 <= (others => '0');
        P_HR_NS726 <= (others => '0');	
			
        P_EDA_NS1 <= (others => '0');
        P_EDA_NS2 <= (others => '0');
        P_EDA_NS3 <= (others => '0');
        P_EDA_NS4 <= (others => '0');
        P_EDA_NS5 <= (others => '0');
        P_EDA_NS6 <= (others => '0');
        P_EDA_NS7 <= (others => '0');
        P_EDA_NS8 <= (others => '0');
        P_EDA_NS9 <= (others => '0');
        P_EDA_NS10 <= (others => '0');
        P_EDA_NS11 <= (others => '0');
        P_EDA_NS12 <= (others => '0');
        P_EDA_NS13 <= (others => '0');
        P_EDA_NS14 <= (others => '0');
        P_EDA_NS15 <= (others => '0');
        P_EDA_NS16 <= (others => '0');
        P_EDA_NS17 <= (others => '0');
        P_EDA_NS18 <= (others => '0');
        P_EDA_NS19 <= (others => '0');
        P_EDA_NS20 <= (others => '0');
        P_EDA_NS21 <= (others => '0');
        P_EDA_NS22 <= (others => '0');
        P_EDA_NS23 <= (others => '0');
        P_EDA_NS24 <= (others => '0');
        P_EDA_NS25 <= (others => '0');
        P_EDA_NS26 <= (others => '0');
        P_EDA_NS27 <= (others => '0');
        P_EDA_NS28 <= (others => '0');
        P_EDA_NS29 <= (others => '0');
        P_EDA_NS30 <= (others => '0');
        P_EDA_NS31 <= (others => '0');
        P_EDA_NS32 <= (others => '0');
        P_EDA_NS33 <= (others => '0');
        P_EDA_NS34 <= (others => '0');
        P_EDA_NS35 <= (others => '0');
        P_EDA_NS36 <= (others => '0');
        P_EDA_NS37 <= (others => '0');
        P_EDA_NS38 <= (others => '0');
        P_EDA_NS39 <= (others => '0');
        P_EDA_NS40 <= (others => '0');
        P_EDA_NS41 <= (others => '0');
        P_EDA_NS42 <= (others => '0');
        P_EDA_NS43 <= (others => '0');
        P_EDA_NS44 <= (others => '0');
        P_EDA_NS45 <= (others => '0');
        P_EDA_NS46 <= (others => '0');
        P_EDA_NS47 <= (others => '0');
        P_EDA_NS48 <= (others => '0');
        P_EDA_NS49 <= (others => '0');
        P_EDA_NS50 <= (others => '0');
        P_EDA_NS51 <= (others => '0');
        P_EDA_NS52 <= (others => '0');
        P_EDA_NS53 <= (others => '0');
        P_EDA_NS54 <= (others => '0');
        P_EDA_NS55 <= (others => '0');
        P_EDA_NS56 <= (others => '0');
        P_EDA_NS57 <= (others => '0');
        P_EDA_NS58 <= (others => '0');
        P_EDA_NS59 <= (others => '0');
        P_EDA_NS60 <= (others => '0');
        P_EDA_NS61 <= (others => '0');
        P_EDA_NS62 <= (others => '0');
        P_EDA_NS63 <= (others => '0');
        P_EDA_NS64 <= (others => '0');
        P_EDA_NS65 <= (others => '0');
        P_EDA_NS66 <= (others => '0');
        P_EDA_NS67 <= (others => '0');
        P_EDA_NS68 <= (others => '0');
        P_EDA_NS69 <= (others => '0');
        P_EDA_NS70 <= (others => '0');
        P_EDA_NS71 <= (others => '0');
        P_EDA_NS72 <= (others => '0');
        P_EDA_NS73 <= (others => '0');
        P_EDA_NS74 <= (others => '0');
        P_EDA_NS75 <= (others => '0');
        P_EDA_NS76 <= (others => '0');
        P_EDA_NS77 <= (others => '0');
        P_EDA_NS78 <= (others => '0');
        P_EDA_NS79 <= (others => '0');
        P_EDA_NS80 <= (others => '0');
        P_EDA_NS81 <= (others => '0');
        P_EDA_NS82 <= (others => '0');
        P_EDA_NS83 <= (others => '0');
        P_EDA_NS84 <= (others => '0');
        P_EDA_NS85 <= (others => '0');
        P_EDA_NS86 <= (others => '0');
        P_EDA_NS87 <= (others => '0');
        P_EDA_NS88 <= (others => '0');
        P_EDA_NS89 <= (others => '0');
        P_EDA_NS90 <= (others => '0');
        P_EDA_NS91 <= (others => '0');
        P_EDA_NS92 <= (others => '0');
        P_EDA_NS93 <= (others => '0');
        P_EDA_NS94 <= (others => '0');
        P_EDA_NS95 <= (others => '0');
        P_EDA_NS96 <= (others => '0');
        P_EDA_NS97 <= (others => '0');
        P_EDA_NS98 <= (others => '0');
        P_EDA_NS99 <= (others => '0');
        P_EDA_NS100 <= (others => '0');
        P_EDA_NS101 <= (others => '0');
        P_EDA_NS102 <= (others => '0');
        P_EDA_NS103 <= (others => '0');
        P_EDA_NS104 <= (others => '0');
        P_EDA_NS105 <= (others => '0');
        P_EDA_NS106 <= (others => '0');
        P_EDA_NS107 <= (others => '0');
        P_EDA_NS108 <= (others => '0');
        P_EDA_NS109 <= (others => '0');
        P_EDA_NS110 <= (others => '0');

		P_TEMP_NS <= (others => '0');	
		P_EDA_NS <= (others => '0');	
		P_HR_NS <= (others => '0');		
		
		not_stress_score <= (others => '0');		
			
		elsif (rising_edge(clk)) then
		if state = NORMAL then
			case temp is
				when "011100000" => P_TEMP_NS <= "0000000001" + P_TEMP_NS1;
				when "011100001" => P_TEMP_NS <= "0000001000" + P_TEMP_NS2;
				when "011100010" => P_TEMP_NS <= "0000100001" + P_TEMP_NS3;
				when "011100011" => P_TEMP_NS <= "0001010100" + P_TEMP_NS4;
				when "011100100" => P_TEMP_NS <= "0001000110" + P_TEMP_NS5;
				when "011100101" => P_TEMP_NS <= "0000010100" + P_TEMP_NS6;
				when "011100110" => P_TEMP_NS <= "0000011010" + P_TEMP_NS7;
				when "011100111" => P_TEMP_NS <= "0000010010" + P_TEMP_NS8;
				when "011101000" => P_TEMP_NS <= "0000000110" + P_TEMP_NS9;
				when "011101001" => P_TEMP_NS <= "0000001010" + P_TEMP_NS10;
				when "011101010" => P_TEMP_NS <= "0000000110" + P_TEMP_NS11;
				when "011101011" => P_TEMP_NS <= "0000000001" + P_TEMP_NS12;
				when "011101100" => P_TEMP_NS <= "0000000001" + P_TEMP_NS13;
				when "011101101" => P_TEMP_NS <= "0000000001" + P_TEMP_NS14;
				when "011101110" => P_TEMP_NS <= "0000000010" + P_TEMP_NS15;
				when "011101111" => P_TEMP_NS <= "0000000010" + P_TEMP_NS16;
				when "011110000" => P_TEMP_NS <= "0000000010" + P_TEMP_NS17;
				when "011110001" => P_TEMP_NS <= "0000000010" + P_TEMP_NS18;
				when "011110010" => P_TEMP_NS <= "0000000010" + P_TEMP_NS19;
				when "011110011" => P_TEMP_NS <= "0000000010" + P_TEMP_NS20;
				when "011110100" => P_TEMP_NS <= "0000000010" + P_TEMP_NS21;
				when "011110101" => P_TEMP_NS <= "0000000010" + P_TEMP_NS22;
				when "011110110" => P_TEMP_NS <= "0000001101" + P_TEMP_NS23;
				when "011110111" => P_TEMP_NS <= "0000111000" + P_TEMP_NS24;
				when "011111000" => P_TEMP_NS <= "0000101101" + P_TEMP_NS25;
				when "011111001" => P_TEMP_NS <= "0000010011" + P_TEMP_NS26;
				when "011111010" => P_TEMP_NS <= "0000101000" + P_TEMP_NS27;
				when "011111011" => P_TEMP_NS <= "0001111011" + P_TEMP_NS28;
				when "011111100" => P_TEMP_NS <= "0000101001" + P_TEMP_NS29;
				when "011111101" => P_TEMP_NS <= "0000111011" + P_TEMP_NS30;
				when "011111110" => P_TEMP_NS <= "0000100000" + P_TEMP_NS31;
				when "011111111" => P_TEMP_NS <= "0000100110" + P_TEMP_NS32;
				when "100000000" => P_TEMP_NS <= "0001001111" + P_TEMP_NS33;
				when "100000001" => P_TEMP_NS <= "0001000110" + P_TEMP_NS34;
				when "100000010" => P_TEMP_NS <= "0000010101" + P_TEMP_NS35;
				when "100000011" => P_TEMP_NS <= "0000001111" + P_TEMP_NS36;
				when "100000100" => P_TEMP_NS <= "0000010100" + P_TEMP_NS37;
				when "100000101" => P_TEMP_NS <= "0000110110" + P_TEMP_NS38;
				when "100000110" => P_TEMP_NS <= "0010100101" + P_TEMP_NS39;
				when "100000111" => P_TEMP_NS <= "0011001000" + P_TEMP_NS40;
				when "100001000" => P_TEMP_NS <= "0011100001" + P_TEMP_NS41;
				when "100001001" => P_TEMP_NS <= "0010110110" + P_TEMP_NS42;
				when "100001010" => P_TEMP_NS <= "0011111000" + P_TEMP_NS43;
				when "100001011" => P_TEMP_NS <= "0011100110" + P_TEMP_NS44;
				when "100001100" => P_TEMP_NS <= "0110100010" + P_TEMP_NS45;
				when "100001101" => P_TEMP_NS <= "0111101001" + P_TEMP_NS46;
				when "100001110" => P_TEMP_NS <= "1000001111" + P_TEMP_NS47;
				when "100001111" => P_TEMP_NS <= "1000010110" + P_TEMP_NS48;
				when "100010000" => P_TEMP_NS <= "1001001101" + P_TEMP_NS49;
				when "100010001" => P_TEMP_NS <= "1001100001" + P_TEMP_NS50;
				when "100010010" => P_TEMP_NS <= "1011011010" + P_TEMP_NS51;
				when "100010011" => P_TEMP_NS <= "1011000110" + P_TEMP_NS52;
				when "100010100" => P_TEMP_NS <= "1001011001" + P_TEMP_NS53;
				when "100010101" => P_TEMP_NS <= "0111101001" + P_TEMP_NS54;
				when "100010110" => P_TEMP_NS <= "1000000011" + P_TEMP_NS55;
				when "100010111" => P_TEMP_NS <= "1000001010" + P_TEMP_NS56;
				when "100011000" => P_TEMP_NS <= "1011111001" + P_TEMP_NS57;
				when "100011001" => P_TEMP_NS <= "0001100110" + P_TEMP_NS58;
				when "100011010" => P_TEMP_NS <= "0000001101" + P_TEMP_NS59;
				when "100011011" => P_TEMP_NS <= "0000100110" + P_TEMP_NS60;
				when "100011100" => P_TEMP_NS <= "0000111100" + P_TEMP_NS61;
				when "100011101" => P_TEMP_NS <= "0000010001" + P_TEMP_NS62;
				when "100011110" => P_TEMP_NS <= "0000000001" + P_TEMP_NS63;
				when  others     => P_TEMP_NS <= "000000000001";
			end case;	
		
        case hr is
				when "00000000001" => P_HR_NS <= "0000001" + P_HR_NS1;
				when "00000000011" => P_HR_NS <= "0000001" + P_HR_NS2;
				when "00000000100" => P_HR_NS <= "0000001" + P_HR_NS3;
				when "00000000111" => P_HR_NS <= "0000001" + P_HR_NS4;
				when "00000001000" => P_HR_NS <= "0000001" + P_HR_NS5;
				when "00000001001" => P_HR_NS <= "0000010" + P_HR_NS6;
				when "00000001010" => P_HR_NS <= "0000001" + P_HR_NS7;
				when "00000001100" => P_HR_NS <= "0000001" + P_HR_NS8;
				when "00000001101" => P_HR_NS <= "0000010" + P_HR_NS9;
				when "00000001110" => P_HR_NS <= "0000001" + P_HR_NS10;
				when "00000001111" => P_HR_NS <= "0000001" + P_HR_NS11;
				when "00000010000" => P_HR_NS <= "0000001" + P_HR_NS12;
				when "00000010001" => P_HR_NS <= "0000010" + P_HR_NS13;
				when "00000010010" => P_HR_NS <= "0000001" + P_HR_NS14;
				when "00000010011" => P_HR_NS <= "0000001" + P_HR_NS15;
				when "00000010101" => P_HR_NS <= "0000001" + P_HR_NS16;
				when "00000010110" => P_HR_NS <= "0000001" + P_HR_NS17;
				when "00000011100" => P_HR_NS <= "0000010" + P_HR_NS18;
				when "00000011101" => P_HR_NS <= "0000001" + P_HR_NS19;
				when "00000011110" => P_HR_NS <= "0000001" + P_HR_NS20;
				when "00000011111" => P_HR_NS <= "0000001" + P_HR_NS21;
				when "00000100000" => P_HR_NS <= "0000001" + P_HR_NS22;
				when "00000100010" => P_HR_NS <= "0000001" + P_HR_NS23;
				when "00000100110" => P_HR_NS <= "0000001" + P_HR_NS24;
				when "00000100111" => P_HR_NS <= "0000001" + P_HR_NS25;
				when "00000101000" => P_HR_NS <= "0000001" + P_HR_NS26;
				when "00000101001" => P_HR_NS <= "0000010" + P_HR_NS27;
				when "00000101010" => P_HR_NS <= "0000001" + P_HR_NS28;
				when "00000101011" => P_HR_NS <= "0000001" + P_HR_NS29;
				when "00000110100" => P_HR_NS <= "0000001" + P_HR_NS30;
				when "00000110101" => P_HR_NS <= "0000001" + P_HR_NS31;
				when "00000111000" => P_HR_NS <= "0000010" + P_HR_NS32;
				when "00000111010" => P_HR_NS <= "0000001" + P_HR_NS33;
				when "00000111100" => P_HR_NS <= "0000001" + P_HR_NS34;
				when "00001000001" => P_HR_NS <= "0000001" + P_HR_NS35;
				when "00001000011" => P_HR_NS <= "0000001" + P_HR_NS36;
				when "00001000100" => P_HR_NS <= "0000001" + P_HR_NS37;
				when "00001000110" => P_HR_NS <= "0000001" + P_HR_NS38;
				when "00001001000" => P_HR_NS <= "0000001" + P_HR_NS39;
				when "00001001100" => P_HR_NS <= "0000001" + P_HR_NS40;
				when "00001001101" => P_HR_NS <= "0000001" + P_HR_NS41;
				when "00001001110" => P_HR_NS <= "0000001" + P_HR_NS42;
				when "00001001111" => P_HR_NS <= "0000001" + P_HR_NS43;
				when "00001010011" => P_HR_NS <= "0000001" + P_HR_NS44;
				when "00001010101" => P_HR_NS <= "0000001" + P_HR_NS45;
				when "00001010110" => P_HR_NS <= "0000001" + P_HR_NS46;
				when "00001011000" => P_HR_NS <= "0000010" + P_HR_NS47;
				when "00001011001" => P_HR_NS <= "0000001" + P_HR_NS48;
				when "00001011010" => P_HR_NS <= "0000001" + P_HR_NS49;
				when "00001011100" => P_HR_NS <= "0000001" + P_HR_NS50;
				when "00001011111" => P_HR_NS <= "0000001" + P_HR_NS51;
				when "00001100000" => P_HR_NS <= "0000001" + P_HR_NS52;
				when "00001100001" => P_HR_NS <= "0000001" + P_HR_NS53;
				when "00001100101" => P_HR_NS <= "0000001" + P_HR_NS54;
				when "00001101000" => P_HR_NS <= "0000001" + P_HR_NS55;
				when "00001101001" => P_HR_NS <= "0000001" + P_HR_NS56;
				when "00001101011" => P_HR_NS <= "0000001" + P_HR_NS57;
				when "00001101100" => P_HR_NS <= "0000001" + P_HR_NS58;
				when "00001101110" => P_HR_NS <= "0000001" + P_HR_NS59;
				when "00001101111" => P_HR_NS <= "0000001" + P_HR_NS60;
				when "00001110000" => P_HR_NS <= "0000001" + P_HR_NS61;
				when "00001110001" => P_HR_NS <= "0000001" + P_HR_NS62;
				when "00001110010" => P_HR_NS <= "0000001" + P_HR_NS63;
				when "00001110101" => P_HR_NS <= "0000001" + P_HR_NS64;
				when "00001110110" => P_HR_NS <= "0000001" + P_HR_NS65;
				when "00001111000" => P_HR_NS <= "0000001" + P_HR_NS66;
				when "00001111011" => P_HR_NS <= "0000001" + P_HR_NS67;
				when "00001111110" => P_HR_NS <= "0000001" + P_HR_NS68;
				when "00001111111" => P_HR_NS <= "0000001" + P_HR_NS69;
				when "00010000000" => P_HR_NS <= "0000001" + P_HR_NS70;
				when "00010000010" => P_HR_NS <= "0000001" + P_HR_NS71;
				when "00010000100" => P_HR_NS <= "0000001" + P_HR_NS72;
				when "00010000101" => P_HR_NS <= "0000001" + P_HR_NS73;
				when "00010000110" => P_HR_NS <= "0000001" + P_HR_NS74;
				when "00010000111" => P_HR_NS <= "0000001" + P_HR_NS75;
				when "00010001001" => P_HR_NS <= "0000001" + P_HR_NS76;
				when "00010001010" => P_HR_NS <= "0000001" + P_HR_NS77;
				when "00010001011" => P_HR_NS <= "0000001" + P_HR_NS78;
				when "00010001100" => P_HR_NS <= "0000010" + P_HR_NS79;
				when "00010001101" => P_HR_NS <= "0000001" + P_HR_NS80;
				when "00010001111" => P_HR_NS <= "0000001" + P_HR_NS81;
				when "00010010000" => P_HR_NS <= "0000001" + P_HR_NS82;
				when "00010010001" => P_HR_NS <= "0000001" + P_HR_NS83;
				when "00010010010" => P_HR_NS <= "0000001" + P_HR_NS84;
				when "00010010011" => P_HR_NS <= "0000001" + P_HR_NS85;
				when "00010010100" => P_HR_NS <= "0000010" + P_HR_NS86;
				when "00010010101" => P_HR_NS <= "0000001" + P_HR_NS87;
				when "00010010110" => P_HR_NS <= "0000001" + P_HR_NS88;
				when "00010010111" => P_HR_NS <= "0000001" + P_HR_NS89;
				when "00010011001" => P_HR_NS <= "0000001" + P_HR_NS90;
				when "00010011100" => P_HR_NS <= "0000001" + P_HR_NS91;
				when "00010011110" => P_HR_NS <= "0000001" + P_HR_NS92;
				when "00010011111" => P_HR_NS <= "0000001" + P_HR_NS93;
				when "00010100001" => P_HR_NS <= "0000010" + P_HR_NS94;
				when "00010100010" => P_HR_NS <= "0000001" + P_HR_NS95;
				when "00010100011" => P_HR_NS <= "0000001" + P_HR_NS96;
				when "00010100100" => P_HR_NS <= "0000001" + P_HR_NS97;
				when "00010100101" => P_HR_NS <= "0000010" + P_HR_NS98;
				when "00010100110" => P_HR_NS <= "0000010" + P_HR_NS99;
				when "00010100111" => P_HR_NS <= "0000001" + P_HR_NS100;
				when "00010101000" => P_HR_NS <= "0000010" + P_HR_NS101;
				when "00010101001" => P_HR_NS <= "0000010" + P_HR_NS102;
				when "00010101010" => P_HR_NS <= "0000010" + P_HR_NS103;
				when "00010101011" => P_HR_NS <= "0000011" + P_HR_NS104;
				when "00010101101" => P_HR_NS <= "0000010" + P_HR_NS105;
				when "00010101110" => P_HR_NS <= "0000010" + P_HR_NS106;
				when "00010101111" => P_HR_NS <= "0000011" + P_HR_NS107;
				when "00010110000" => P_HR_NS <= "0000010" + P_HR_NS108;
				when "00010110001" => P_HR_NS <= "0000010" + P_HR_NS109;
				when "00010110010" => P_HR_NS <= "0000010" + P_HR_NS110;
				when "00010110011" => P_HR_NS <= "0000100" + P_HR_NS111;
				when "00010110100" => P_HR_NS <= "0000010" + P_HR_NS112;
				when "00010110101" => P_HR_NS <= "0000010" + P_HR_NS113;
				when "00010110110" => P_HR_NS <= "0000010" + P_HR_NS114;
				when "00010110111" => P_HR_NS <= "0000010" + P_HR_NS115;
				when "00010111000" => P_HR_NS <= "0000010" + P_HR_NS116;
				when "00010111001" => P_HR_NS <= "0000010" + P_HR_NS117;
				when "00010111010" => P_HR_NS <= "0000010" + P_HR_NS118;
				when "00010111011" => P_HR_NS <= "0000010" + P_HR_NS119;
				when "00010111100" => P_HR_NS <= "0000010" + P_HR_NS120;
				when "00010111101" => P_HR_NS <= "0000001" + P_HR_NS121;
				when "00010111110" => P_HR_NS <= "0000010" + P_HR_NS122;
				when "00010111111" => P_HR_NS <= "0000010" + P_HR_NS123;
				when "00011000000" => P_HR_NS <= "0000001" + P_HR_NS124;
				when "00011000001" => P_HR_NS <= "0000010" + P_HR_NS125;
				when "00011000010" => P_HR_NS <= "0000001" + P_HR_NS126;
				when "00011000011" => P_HR_NS <= "0000010" + P_HR_NS127;
				when "00011000100" => P_HR_NS <= "0000010" + P_HR_NS128;
				when "00011000101" => P_HR_NS <= "0000010" + P_HR_NS129;
				when "00011000110" => P_HR_NS <= "0000001" + P_HR_NS130;
				when "00011000111" => P_HR_NS <= "0000001" + P_HR_NS131;
				when "00011001000" => P_HR_NS <= "0000010" + P_HR_NS132;
				when "00011001001" => P_HR_NS <= "0000001" + P_HR_NS133;
				when "00011001010" => P_HR_NS <= "0000010" + P_HR_NS134;
				when "00011001011" => P_HR_NS <= "0000001" + P_HR_NS135;
				when "00011001100" => P_HR_NS <= "0000010" + P_HR_NS136;
				when "00011001101" => P_HR_NS <= "0000001" + P_HR_NS137;
				when "00011001111" => P_HR_NS <= "0000010" + P_HR_NS138;
				when "00011010000" => P_HR_NS <= "0000010" + P_HR_NS139;
				when "00011010001" => P_HR_NS <= "0000001" + P_HR_NS140;
				when "00011010010" => P_HR_NS <= "0000001" + P_HR_NS141;
				when "00011010011" => P_HR_NS <= "0000001" + P_HR_NS142;
				when "00011010100" => P_HR_NS <= "0000010" + P_HR_NS143;
				when "00011010101" => P_HR_NS <= "0000010" + P_HR_NS144;
				when "00011010110" => P_HR_NS <= "0000001" + P_HR_NS145;
				when "00011010111" => P_HR_NS <= "0000001" + P_HR_NS146;
				when "00011011000" => P_HR_NS <= "0000001" + P_HR_NS147;
				when "00011011001" => P_HR_NS <= "0000001" + P_HR_NS148;
				when "00011011011" => P_HR_NS <= "0000001" + P_HR_NS149;
				when "00011100000" => P_HR_NS <= "0000001" + P_HR_NS150;
				when "00011100010" => P_HR_NS <= "0000010" + P_HR_NS151;
				when "00011100011" => P_HR_NS <= "0000001" + P_HR_NS152;
				when "00011100100" => P_HR_NS <= "0000001" + P_HR_NS153;
				when "00011100101" => P_HR_NS <= "0000001" + P_HR_NS154;
				when "00011100110" => P_HR_NS <= "0000001" + P_HR_NS155;
				when "00011100111" => P_HR_NS <= "0000001" + P_HR_NS156;
				when "00011101000" => P_HR_NS <= "0000001" + P_HR_NS157;
				when "00011101001" => P_HR_NS <= "0000001" + P_HR_NS158;
				when "00011101010" => P_HR_NS <= "0000001" + P_HR_NS159;
				when "00011101011" => P_HR_NS <= "0000001" + P_HR_NS160;
				when "00011101101" => P_HR_NS <= "0000001" + P_HR_NS161;
				when "00011101111" => P_HR_NS <= "0000001" + P_HR_NS162;
				when "00011110000" => P_HR_NS <= "0000010" + P_HR_NS163;
				when "00011110011" => P_HR_NS <= "0000001" + P_HR_NS164;
				when "00011110101" => P_HR_NS <= "0000001" + P_HR_NS165;
				when "00011110110" => P_HR_NS <= "0000001" + P_HR_NS166;
				when "00011111000" => P_HR_NS <= "0000001" + P_HR_NS167;
				when "00011111001" => P_HR_NS <= "0000010" + P_HR_NS168;
				when "00011111010" => P_HR_NS <= "0000001" + P_HR_NS169;
				when "00011111011" => P_HR_NS <= "0000010" + P_HR_NS170;
				when "00011111100" => P_HR_NS <= "0000001" + P_HR_NS171;
				when "00011111101" => P_HR_NS <= "0000010" + P_HR_NS172;
				when "00011111110" => P_HR_NS <= "0000001" + P_HR_NS173;
				when "00011111111" => P_HR_NS <= "0000001" + P_HR_NS174;
				when "00100000000" => P_HR_NS <= "0000010" + P_HR_NS175;
				when "00100000001" => P_HR_NS <= "0000010" + P_HR_NS176;
				when "00100000010" => P_HR_NS <= "0000010" + P_HR_NS177;
				when "00100000011" => P_HR_NS <= "0000010" + P_HR_NS178;
				when "00100000100" => P_HR_NS <= "0000011" + P_HR_NS179;
				when "00100000101" => P_HR_NS <= "0000010" + P_HR_NS180;
				when "00100000110" => P_HR_NS <= "0000010" + P_HR_NS181;
				when "00100000111" => P_HR_NS <= "0000001" + P_HR_NS182;
				when "00100001000" => P_HR_NS <= "0000001" + P_HR_NS183;
				when "00100001001" => P_HR_NS <= "0000001" + P_HR_NS184;
				when "00100001010" => P_HR_NS <= "0000011" + P_HR_NS185;
				when "00100001011" => P_HR_NS <= "0000010" + P_HR_NS186;
				when "00100001100" => P_HR_NS <= "0000010" + P_HR_NS187;
				when "00100001101" => P_HR_NS <= "0000011" + P_HR_NS188;
				when "00100001110" => P_HR_NS <= "0000001" + P_HR_NS189;
				when "00100001111" => P_HR_NS <= "0000011" + P_HR_NS190;
				when "00100010000" => P_HR_NS <= "0000010" + P_HR_NS191;
				when "00100010001" => P_HR_NS <= "0000010" + P_HR_NS192;
				when "00100010010" => P_HR_NS <= "0000010" + P_HR_NS193;
				when "00100010011" => P_HR_NS <= "0000001" + P_HR_NS194;
				when "00100010100" => P_HR_NS <= "0000010" + P_HR_NS195;
				when "00100010101" => P_HR_NS <= "0000010" + P_HR_NS196;
				when "00100010110" => P_HR_NS <= "0000010" + P_HR_NS197;
				when "00100010111" => P_HR_NS <= "0000010" + P_HR_NS198;
				when "00100011000" => P_HR_NS <= "0000010" + P_HR_NS199;
				when "00100011001" => P_HR_NS <= "0000010" + P_HR_NS200;
				when "00100011010" => P_HR_NS <= "0000001" + P_HR_NS201;
				when "00100011011" => P_HR_NS <= "0000001" + P_HR_NS202;
				when "00100011100" => P_HR_NS <= "0000001" + P_HR_NS203;
				when "00100011101" => P_HR_NS <= "0000001" + P_HR_NS204;
				when "00100011110" => P_HR_NS <= "0000001" + P_HR_NS205;
				when "00100011111" => P_HR_NS <= "0000001" + P_HR_NS206;
				when "00100100000" => P_HR_NS <= "0000001" + P_HR_NS207;
				when "00100100001" => P_HR_NS <= "0000010" + P_HR_NS208;
				when "00100100010" => P_HR_NS <= "0000001" + P_HR_NS209;
				when "00100100011" => P_HR_NS <= "0000001" + P_HR_NS210;
				when "00100100100" => P_HR_NS <= "0000001" + P_HR_NS211;
				when "00100100101" => P_HR_NS <= "0000001" + P_HR_NS212;
				when "00100100110" => P_HR_NS <= "0000001" + P_HR_NS213;
				when "00100101001" => P_HR_NS <= "0000010" + P_HR_NS214;
				when "00100101010" => P_HR_NS <= "0000001" + P_HR_NS215;
				when "00100101011" => P_HR_NS <= "0000010" + P_HR_NS216;
				when "00100101100" => P_HR_NS <= "0000001" + P_HR_NS217;
				when "00100101101" => P_HR_NS <= "0000001" + P_HR_NS218;
				when "00100101110" => P_HR_NS <= "0000001" + P_HR_NS219;
				when "00100110000" => P_HR_NS <= "0000001" + P_HR_NS220;
				when "00100110010" => P_HR_NS <= "0000001" + P_HR_NS221;
				when "00100110011" => P_HR_NS <= "0000001" + P_HR_NS222;
				when "00100110100" => P_HR_NS <= "0000001" + P_HR_NS223;
				when "00100110110" => P_HR_NS <= "0000001" + P_HR_NS224;
				when "00100111000" => P_HR_NS <= "0000001" + P_HR_NS225;
				when "00100111010" => P_HR_NS <= "0000001" + P_HR_NS226;
				when "00100111011" => P_HR_NS <= "0000010" + P_HR_NS227;
				when "00100111100" => P_HR_NS <= "0000001" + P_HR_NS228;
				when "00100111110" => P_HR_NS <= "0000001" + P_HR_NS229;
				when "00100111111" => P_HR_NS <= "0000001" + P_HR_NS230;
				when "00101000000" => P_HR_NS <= "0000010" + P_HR_NS231;
				when "00101000010" => P_HR_NS <= "0000001" + P_HR_NS232;
				when "00101000011" => P_HR_NS <= "0000001" + P_HR_NS233;
				when "00101000100" => P_HR_NS <= "0000001" + P_HR_NS234;
				when "00101000101" => P_HR_NS <= "0000001" + P_HR_NS235;
				when "00101000110" => P_HR_NS <= "0000001" + P_HR_NS236;
				when "00101000111" => P_HR_NS <= "0000001" + P_HR_NS237;
				when "00101001000" => P_HR_NS <= "0000001" + P_HR_NS238;
				when "00101001011" => P_HR_NS <= "0000010" + P_HR_NS239;
				when "00101001100" => P_HR_NS <= "0000001" + P_HR_NS240;
				when "00101001110" => P_HR_NS <= "0000001" + P_HR_NS241;
				when "00101001111" => P_HR_NS <= "0000001" + P_HR_NS242;
				when "00101010000" => P_HR_NS <= "0000001" + P_HR_NS243;
				when "00101010001" => P_HR_NS <= "0000010" + P_HR_NS244;
				when "00101010010" => P_HR_NS <= "0000010" + P_HR_NS245;
				when "00101010011" => P_HR_NS <= "0000001" + P_HR_NS246;
				when "00101010100" => P_HR_NS <= "0000010" + P_HR_NS247;
				when "00101010101" => P_HR_NS <= "0000001" + P_HR_NS248;
				when "00101010110" => P_HR_NS <= "0000001" + P_HR_NS249;
				when "00101010111" => P_HR_NS <= "0000010" + P_HR_NS250;
				when "00101011000" => P_HR_NS <= "0000010" + P_HR_NS251;
				when "00101011001" => P_HR_NS <= "0000001" + P_HR_NS252;
				when "00101011010" => P_HR_NS <= "0000010" + P_HR_NS253;
				when "00101011011" => P_HR_NS <= "0000010" + P_HR_NS254;
				when "00101011100" => P_HR_NS <= "0000010" + P_HR_NS255;
				when "00101011101" => P_HR_NS <= "0000011" + P_HR_NS256;
				when "00101011110" => P_HR_NS <= "0000010" + P_HR_NS257;
				when "00101011111" => P_HR_NS <= "0000001" + P_HR_NS258;
				when "00101100000" => P_HR_NS <= "0000001" + P_HR_NS259;
				when "00101100001" => P_HR_NS <= "0000010" + P_HR_NS260;
				when "00101100010" => P_HR_NS <= "0000011" + P_HR_NS261;
				when "00101100011" => P_HR_NS <= "0000010" + P_HR_NS262;
				when "00101100100" => P_HR_NS <= "0000010" + P_HR_NS263;
				when "00101100101" => P_HR_NS <= "0000011" + P_HR_NS264;
				when "00101100110" => P_HR_NS <= "0000001" + P_HR_NS265;
				when "00101100111" => P_HR_NS <= "0000100" + P_HR_NS266;
				when "00101101000" => P_HR_NS <= "0000011" + P_HR_NS267;
				when "00101101001" => P_HR_NS <= "0000100" + P_HR_NS268;
				when "00101101010" => P_HR_NS <= "0000100" + P_HR_NS269;
				when "00101101011" => P_HR_NS <= "0000011" + P_HR_NS270;
				when "00101101100" => P_HR_NS <= "0000011" + P_HR_NS271;
				when "00101101101" => P_HR_NS <= "0000011" + P_HR_NS272;
				when "00101101110" => P_HR_NS <= "0000110" + P_HR_NS273;
				when "00101101111" => P_HR_NS <= "0000011" + P_HR_NS274;
				when "00101110000" => P_HR_NS <= "0000101" + P_HR_NS275;
				when "00101110001" => P_HR_NS <= "0000011" + P_HR_NS276;
				when "00101110010" => P_HR_NS <= "0000110" + P_HR_NS277;
				when "00101110011" => P_HR_NS <= "0000011" + P_HR_NS278;
				when "00101110100" => P_HR_NS <= "0000010" + P_HR_NS279;
				when "00101110101" => P_HR_NS <= "0000100" + P_HR_NS280;
				when "00101110110" => P_HR_NS <= "0000100" + P_HR_NS281;
				when "00101110111" => P_HR_NS <= "0000110" + P_HR_NS282;
				when "00101111000" => P_HR_NS <= "0000101" + P_HR_NS283;
				when "00101111001" => P_HR_NS <= "0000100" + P_HR_NS284;
				when "00101111010" => P_HR_NS <= "0000101" + P_HR_NS285;
				when "00101111011" => P_HR_NS <= "0000011" + P_HR_NS286;
				when "00101111100" => P_HR_NS <= "0000011" + P_HR_NS287;
				when "00101111101" => P_HR_NS <= "0001000" + P_HR_NS288;
				when "00101111110" => P_HR_NS <= "0000100" + P_HR_NS289;
				when "00101111111" => P_HR_NS <= "0000011" + P_HR_NS290;
				when "00110000000" => P_HR_NS <= "0000110" + P_HR_NS291;
				when "00110000001" => P_HR_NS <= "0000100" + P_HR_NS292;
				when "00110000010" => P_HR_NS <= "0000011" + P_HR_NS293;
				when "00110000011" => P_HR_NS <= "0000110" + P_HR_NS294;
				when "00110000100" => P_HR_NS <= "0001000" + P_HR_NS295;
				when "00110000101" => P_HR_NS <= "0000100" + P_HR_NS296;
				when "00110000110" => P_HR_NS <= "0000110" + P_HR_NS297;
				when "00110000111" => P_HR_NS <= "0000110" + P_HR_NS298;
				when "00110001000" => P_HR_NS <= "0000101" + P_HR_NS299;
				when "00110001001" => P_HR_NS <= "0001011" + P_HR_NS300;
				when "00110001010" => P_HR_NS <= "0000110" + P_HR_NS301;
				when "00110001011" => P_HR_NS <= "0000110" + P_HR_NS302;
				when "00110001100" => P_HR_NS <= "0000111" + P_HR_NS303;
				when "00110001101" => P_HR_NS <= "0000110" + P_HR_NS304;
				when "00110001110" => P_HR_NS <= "0001001" + P_HR_NS305;
				when "00110001111" => P_HR_NS <= "0000101" + P_HR_NS306;
				when "00110010000" => P_HR_NS <= "0001011" + P_HR_NS307;
				when "00110010001" => P_HR_NS <= "0001000" + P_HR_NS308;
				when "00110010010" => P_HR_NS <= "0001001" + P_HR_NS309;
				when "00110010011" => P_HR_NS <= "0001011" + P_HR_NS310;
				when "00110010100" => P_HR_NS <= "0001001" + P_HR_NS311;
				when "00110010101" => P_HR_NS <= "0001001" + P_HR_NS312;
				when "00110010110" => P_HR_NS <= "0001000" + P_HR_NS313;
				when "00110010111" => P_HR_NS <= "0001011" + P_HR_NS314;
				when "00110011000" => P_HR_NS <= "0000111" + P_HR_NS315;
				when "00110011001" => P_HR_NS <= "0001010" + P_HR_NS316;
				when "00110011010" => P_HR_NS <= "0001010" + P_HR_NS317;
				when "00110011011" => P_HR_NS <= "0001000" + P_HR_NS318;
				when "00110011100" => P_HR_NS <= "0001000" + P_HR_NS319;
				when "00110011101" => P_HR_NS <= "0001010" + P_HR_NS320;
				when "00110011110" => P_HR_NS <= "0001001" + P_HR_NS321;
				when "00110011111" => P_HR_NS <= "0001001" + P_HR_NS322;
				when "00110100000" => P_HR_NS <= "0001010" + P_HR_NS323;
				when "00110100001" => P_HR_NS <= "0001001" + P_HR_NS324;
				when "00110100010" => P_HR_NS <= "0001010" + P_HR_NS325;
				when "00110100011" => P_HR_NS <= "0001010" + P_HR_NS326;
				when "00110100100" => P_HR_NS <= "0000101" + P_HR_NS327;
				when "00110100101" => P_HR_NS <= "0001100" + P_HR_NS328;
				when "00110100110" => P_HR_NS <= "0001100" + P_HR_NS329;
				when "00110100111" => P_HR_NS <= "0001010" + P_HR_NS330;
				when "00110101000" => P_HR_NS <= "0001011" + P_HR_NS331;
				when "00110101001" => P_HR_NS <= "0001011" + P_HR_NS332;
				when "00110101010" => P_HR_NS <= "0001110" + P_HR_NS333;
				when "00110101011" => P_HR_NS <= "0001100" + P_HR_NS334;
				when "00110101100" => P_HR_NS <= "0000111" + P_HR_NS335;
				when "00110101101" => P_HR_NS <= "0001111" + P_HR_NS336;
				when "00110101110" => P_HR_NS <= "0001101" + P_HR_NS337;
				when "00110101111" => P_HR_NS <= "0001000" + P_HR_NS338;
				when "00110110000" => P_HR_NS <= "0001111" + P_HR_NS339;
				when "00110110001" => P_HR_NS <= "0000101" + P_HR_NS340;
				when "00110110010" => P_HR_NS <= "0001111" + P_HR_NS341;
				when "00110110011" => P_HR_NS <= "0001110" + P_HR_NS342;
				when "00110110100" => P_HR_NS <= "0010001" + P_HR_NS343;
				when "00110110101" => P_HR_NS <= "0001010" + P_HR_NS344;
				when "00110110110" => P_HR_NS <= "0010000" + P_HR_NS345;
				when "00110110111" => P_HR_NS <= "0010000" + P_HR_NS346;
				when "00110111000" => P_HR_NS <= "0001111" + P_HR_NS347;
				when "00110111001" => P_HR_NS <= "0001001" + P_HR_NS348;
				when "00110111010" => P_HR_NS <= "0001101" + P_HR_NS349;
				when "00110111011" => P_HR_NS <= "0010001" + P_HR_NS350;
				when "00110111100" => P_HR_NS <= "0010011" + P_HR_NS351;
				when "00110111101" => P_HR_NS <= "0001001" + P_HR_NS352;
				when "00110111110" => P_HR_NS <= "0010001" + P_HR_NS353;
				when "00110111111" => P_HR_NS <= "0010001" + P_HR_NS354;
				when "00111000000" => P_HR_NS <= "0001011" + P_HR_NS355;
				when "00111000001" => P_HR_NS <= "0010100" + P_HR_NS356;
				when "00111000010" => P_HR_NS <= "0010001" + P_HR_NS357;
				when "00111000011" => P_HR_NS <= "0001011" + P_HR_NS358;
				when "00111000100" => P_HR_NS <= "0010101" + P_HR_NS359;
				when "00111000101" => P_HR_NS <= "0010111" + P_HR_NS360;
				when "00111000110" => P_HR_NS <= "0001011" + P_HR_NS361;
				when "00111000111" => P_HR_NS <= "0010111" + P_HR_NS362;
				when "00111001000" => P_HR_NS <= "0001011" + P_HR_NS363;
				when "00111001001" => P_HR_NS <= "0011000" + P_HR_NS364;
				when "00111001010" => P_HR_NS <= "0010111" + P_HR_NS365;
				when "00111001011" => P_HR_NS <= "0001001" + P_HR_NS366;
				when "00111001100" => P_HR_NS <= "0011010" + P_HR_NS367;
				when "00111001101" => P_HR_NS <= "0001011" + P_HR_NS368;
				when "00111001110" => P_HR_NS <= "0011100" + P_HR_NS369;
				when "00111001111" => P_HR_NS <= "0011100" + P_HR_NS370;
				when "00111010000" => P_HR_NS <= "0001101" + P_HR_NS371;
				when "00111010001" => P_HR_NS <= "0011000" + P_HR_NS372;
				when "00111010010" => P_HR_NS <= "0001101" + P_HR_NS373;
				when "00111010011" => P_HR_NS <= "0011111" + P_HR_NS374;
				when "00111010100" => P_HR_NS <= "0001110" + P_HR_NS375;
				when "00111010101" => P_HR_NS <= "0011110" + P_HR_NS376;
				when "00111010110" => P_HR_NS <= "0001110" + P_HR_NS377;
				when "00111010111" => P_HR_NS <= "0011100" + P_HR_NS378;
				when "00111011000" => P_HR_NS <= "0010001" + P_HR_NS379;
				when "00111011001" => P_HR_NS <= "0100101" + P_HR_NS380;
				when "00111011010" => P_HR_NS <= "0010100" + P_HR_NS381;
				when "00111011011" => P_HR_NS <= "0100000" + P_HR_NS382;
				when "00111011100" => P_HR_NS <= "0010010" + P_HR_NS383;
				when "00111011101" => P_HR_NS <= "0100101" + P_HR_NS384;
				when "00111011110" => P_HR_NS <= "0010101" + P_HR_NS385;
				when "00111011111" => P_HR_NS <= "0100010" + P_HR_NS386;
				when "00111100000" => P_HR_NS <= "0001111" + P_HR_NS387;
				when "00111100001" => P_HR_NS <= "0100110" + P_HR_NS388;
				when "00111100010" => P_HR_NS <= "0010000" + P_HR_NS389;
				when "00111100011" => P_HR_NS <= "0100011" + P_HR_NS390;
				when "00111100100" => P_HR_NS <= "0010000" + P_HR_NS391;
				when "00111100101" => P_HR_NS <= "0010110" + P_HR_NS392;
				when "00111100110" => P_HR_NS <= "0101010" + P_HR_NS393;
				when "00111100111" => P_HR_NS <= "0010000" + P_HR_NS394;
				when "00111101000" => P_HR_NS <= "0101100" + P_HR_NS395;
				when "00111101001" => P_HR_NS <= "0010011" + P_HR_NS396;
				when "00111101010" => P_HR_NS <= "0011000" + P_HR_NS397;
				when "00111101011" => P_HR_NS <= "0110000" + P_HR_NS398;
				when "00111101100" => P_HR_NS <= "0010101" + P_HR_NS399;
				when "00111101101" => P_HR_NS <= "0101111" + P_HR_NS400;
				when "00111101110" => P_HR_NS <= "0011000" + P_HR_NS401;
				when "00111101111" => P_HR_NS <= "0011011" + P_HR_NS402;
				when "00111110000" => P_HR_NS <= "0101110" + P_HR_NS403;
				when "00111110001" => P_HR_NS <= "0010101" + P_HR_NS404;
				when "00111110010" => P_HR_NS <= "0001111" + P_HR_NS405;
				when "00111110011" => P_HR_NS <= "0110001" + P_HR_NS406;
				when "00111110100" => P_HR_NS <= "0011001" + P_HR_NS407;
				when "00111110101" => P_HR_NS <= "0101111" + P_HR_NS408;
				when "00111110110" => P_HR_NS <= "0011110" + P_HR_NS409;
				when "00111110111" => P_HR_NS <= "0011100" + P_HR_NS410;
				when "00111111000" => P_HR_NS <= "0010110" + P_HR_NS411;
				when "00111111001" => P_HR_NS <= "0110111" + P_HR_NS412;
				when "00111111010" => P_HR_NS <= "0011101" + P_HR_NS413;
				when "00111111011" => P_HR_NS <= "0011011" + P_HR_NS414;
				when "00111111100" => P_HR_NS <= "0101100" + P_HR_NS415;
				when "00111111101" => P_HR_NS <= "0010111" + P_HR_NS416;
				when "00111111110" => P_HR_NS <= "0011101" + P_HR_NS417;
				when "00111111111" => P_HR_NS <= "0111000" + P_HR_NS418;
				when "01000000000" => P_HR_NS <= "0011001" + P_HR_NS419;
				when "01000000001" => P_HR_NS <= "0011001" + P_HR_NS420;
				when "01000000010" => P_HR_NS <= "0011111" + P_HR_NS421;
				when "01000000011" => P_HR_NS <= "0111111" + P_HR_NS422;
				when "01000000100" => P_HR_NS <= "0011111" + P_HR_NS423;
				when "01000000101" => P_HR_NS <= "0011100" + P_HR_NS424;
				when "01000000110" => P_HR_NS <= "0011011" + P_HR_NS425;
				when "01000000111" => P_HR_NS <= "0111100" + P_HR_NS426;
				when "01000001000" => P_HR_NS <= "0011011" + P_HR_NS427;
				when "01000001001" => P_HR_NS <= "0011111" + P_HR_NS428;
				when "01000001010" => P_HR_NS <= "0011101" + P_HR_NS429;
				when "01000001011" => P_HR_NS <= "0111110" + P_HR_NS430;
				when "01000001100" => P_HR_NS <= "0011100" + P_HR_NS431;
				when "01000001101" => P_HR_NS <= "0011101" + P_HR_NS432;
				when "01000001110" => P_HR_NS <= "0011101" + P_HR_NS433;
				when "01000001111" => P_HR_NS <= "0111000" + P_HR_NS434;
				when "01000010000" => P_HR_NS <= "0011011" + P_HR_NS435;
				when "01000010001" => P_HR_NS <= "0011011" + P_HR_NS436;
				when "01000010010" => P_HR_NS <= "0011110" + P_HR_NS437;
				when "01000010011" => P_HR_NS <= "0100001" + P_HR_NS438;
				when "01000010100" => P_HR_NS <= "1000100" + P_HR_NS439;
				when "01000010101" => P_HR_NS <= "0100010" + P_HR_NS440;
				when "01000010110" => P_HR_NS <= "0100100" + P_HR_NS441;
				when "01000010111" => P_HR_NS <= "0011111" + P_HR_NS442;
				when "01000011000" => P_HR_NS <= "0100001" + P_HR_NS443;
				when "01000011001" => P_HR_NS <= "0011010" + P_HR_NS444;
				when "01000011010" => P_HR_NS <= "1000010" + P_HR_NS445;
				when "01000011011" => P_HR_NS <= "0100000" + P_HR_NS446;
				when "01000011100" => P_HR_NS <= "0100010" + P_HR_NS447;
				when "01000011101" => P_HR_NS <= "0100000" + P_HR_NS448;
				when "01000011110" => P_HR_NS <= "0100000" + P_HR_NS449;
				when "01000011111" => P_HR_NS <= "0100000" + P_HR_NS450;
				when "01000100000" => P_HR_NS <= "0100001" + P_HR_NS451;
				when "01000100001" => P_HR_NS <= "1000100" + P_HR_NS452;
				when "01000100010" => P_HR_NS <= "0100010" + P_HR_NS453;
				when "01000100011" => P_HR_NS <= "0011111" + P_HR_NS454;
				when "01000100100" => P_HR_NS <= "0100100" + P_HR_NS455;
				when "01000100101" => P_HR_NS <= "0011100" + P_HR_NS456;
				when "01000100110" => P_HR_NS <= "0101000" + P_HR_NS457;
				when "01000100111" => P_HR_NS <= "0100001" + P_HR_NS458;
				when "01000101000" => P_HR_NS <= "0011110" + P_HR_NS459;
				when "01000101001" => P_HR_NS <= "0100000" + P_HR_NS460;
				when "01000101010" => P_HR_NS <= "1000111" + P_HR_NS461;
				when "01000101011" => P_HR_NS <= "0100010" + P_HR_NS462;
				when "01000101100" => P_HR_NS <= "0100110" + P_HR_NS463;
				when "01000101101" => P_HR_NS <= "0100100" + P_HR_NS464;
				when "01000101110" => P_HR_NS <= "0011011" + P_HR_NS465;
				when "01000101111" => P_HR_NS <= "0101000" + P_HR_NS466;
				when "01000110000" => P_HR_NS <= "0100010" + P_HR_NS467;
				when "01000110001" => P_HR_NS <= "0100100" + P_HR_NS468;
				when "01000110010" => P_HR_NS <= "0100111" + P_HR_NS469;
				when "01000110011" => P_HR_NS <= "0100011" + P_HR_NS470;
				when "01000110100" => P_HR_NS <= "0100100" + P_HR_NS471;
				when "01000110101" => P_HR_NS <= "0100010" + P_HR_NS472;
				when "01000110110" => P_HR_NS <= "0100010" + P_HR_NS473;
				when "01000110111" => P_HR_NS <= "0100001" + P_HR_NS474;
				when "01000111000" => P_HR_NS <= "0100010" + P_HR_NS475;
				when "01000111001" => P_HR_NS <= "1000010" + P_HR_NS476;
				when "01000111010" => P_HR_NS <= "0101001" + P_HR_NS477;
				when "01000111011" => P_HR_NS <= "0100101" + P_HR_NS478;
				when "01000111100" => P_HR_NS <= "0100011" + P_HR_NS479;
				when "01000111101" => P_HR_NS <= "0100010" + P_HR_NS480;
				when "01000111110" => P_HR_NS <= "0100001" + P_HR_NS481;
				when "01000111111" => P_HR_NS <= "0100010" + P_HR_NS482;
				when "01001000000" => P_HR_NS <= "0100100" + P_HR_NS483;
				when "01001000001" => P_HR_NS <= "0011110" + P_HR_NS484;
				when "01001000010" => P_HR_NS <= "0100110" + P_HR_NS485;
				when "01001000011" => P_HR_NS <= "0100100" + P_HR_NS486;
				when "01001000100" => P_HR_NS <= "0100100" + P_HR_NS487;
				when "01001000101" => P_HR_NS <= "0100100" + P_HR_NS488;
				when "01001000110" => P_HR_NS <= "0100110" + P_HR_NS489;
				when "01001000111" => P_HR_NS <= "0100011" + P_HR_NS490;
				when "01001001000" => P_HR_NS <= "0011100" + P_HR_NS491;
				when "01001001001" => P_HR_NS <= "0100100" + P_HR_NS492;
				when "01001001010" => P_HR_NS <= "0100011" + P_HR_NS493;
				when "01001001011" => P_HR_NS <= "0100100" + P_HR_NS494;
				when "01001001100" => P_HR_NS <= "0100110" + P_HR_NS495;
				when "01001001101" => P_HR_NS <= "0101000" + P_HR_NS496;
				when "01001001111" => P_HR_NS <= "0100111" + P_HR_NS497;
				when "01001010000" => P_HR_NS <= "0101000" + P_HR_NS498;
				when "01001010001" => P_HR_NS <= "0100100" + P_HR_NS499;
				when "01001010010" => P_HR_NS <= "0010110" + P_HR_NS500;
				when "01001010011" => P_HR_NS <= "0101001" + P_HR_NS501;
				when "01001010100" => P_HR_NS <= "0100010" + P_HR_NS502;
				when "01001010101" => P_HR_NS <= "0100010" + P_HR_NS503;
				when "01001010110" => P_HR_NS <= "0100011" + P_HR_NS504;
				when "01001010111" => P_HR_NS <= "0100001" + P_HR_NS505;
				when "01001011000" => P_HR_NS <= "0100111" + P_HR_NS506;
				when "01001011001" => P_HR_NS <= "0100010" + P_HR_NS507;
				when "01001011010" => P_HR_NS <= "0011110" + P_HR_NS508;
				when "01001011011" => P_HR_NS <= "0011100" + P_HR_NS509;
				when "01001011100" => P_HR_NS <= "0100100" + P_HR_NS510;
				when "01001011101" => P_HR_NS <= "0100100" + P_HR_NS511;
				when "01001011110" => P_HR_NS <= "0100101" + P_HR_NS512;
				when "01001100000" => P_HR_NS <= "0100100" + P_HR_NS513;
				when "01001100001" => P_HR_NS <= "0100101" + P_HR_NS514;
				when "01001100010" => P_HR_NS <= "0100010" + P_HR_NS515;
				when "01001100011" => P_HR_NS <= "0011101" + P_HR_NS516;
				when "01001100100" => P_HR_NS <= "0100111" + P_HR_NS517;
				when "01001100101" => P_HR_NS <= "0100001" + P_HR_NS518;
				when "01001100110" => P_HR_NS <= "0011111" + P_HR_NS519;
				when "01001100111" => P_HR_NS <= "0100011" + P_HR_NS520;
				when "01001101001" => P_HR_NS <= "0011101" + P_HR_NS521;
				when "01001101010" => P_HR_NS <= "0100100" + P_HR_NS522;
				when "01001101011" => P_HR_NS <= "0101101" + P_HR_NS523;
				when "01001101100" => P_HR_NS <= "0100111" + P_HR_NS524;
				when "01001101101" => P_HR_NS <= "0100000" + P_HR_NS525;
				when "01001101110" => P_HR_NS <= "0100000" + P_HR_NS526;
				when "01001101111" => P_HR_NS <= "0101010" + P_HR_NS527;
				when "01001110001" => P_HR_NS <= "0100100" + P_HR_NS528;
				when "01001110010" => P_HR_NS <= "0100010" + P_HR_NS529;
				when "01001110011" => P_HR_NS <= "0101000" + P_HR_NS530;
				when "01001110100" => P_HR_NS <= "0100001" + P_HR_NS531;
				when "01001110101" => P_HR_NS <= "0011111" + P_HR_NS532;
				when "01001110110" => P_HR_NS <= "0100101" + P_HR_NS533;
				when "01001111000" => P_HR_NS <= "0100100" + P_HR_NS534;
				when "01001111001" => P_HR_NS <= "0100000" + P_HR_NS535;
				when "01001111010" => P_HR_NS <= "0100010" + P_HR_NS536;
				when "01001111011" => P_HR_NS <= "0100010" + P_HR_NS537;
				when "01001111100" => P_HR_NS <= "0100010" + P_HR_NS538;
				when "01001111110" => P_HR_NS <= "0100010" + P_HR_NS539;
				when "01001111111" => P_HR_NS <= "0100000" + P_HR_NS540;
				when "01010000000" => P_HR_NS <= "0011101" + P_HR_NS541;
				when "01010000001" => P_HR_NS <= "0100100" + P_HR_NS542;
				when "01010000010" => P_HR_NS <= "0100101" + P_HR_NS543;
				when "01010000100" => P_HR_NS <= "0100000" + P_HR_NS544;
				when "01010000101" => P_HR_NS <= "0011101" + P_HR_NS545;
				when "01010000110" => P_HR_NS <= "0100011" + P_HR_NS546;
				when "01010000111" => P_HR_NS <= "0011110" + P_HR_NS547;
				when "01010001001" => P_HR_NS <= "0011100" + P_HR_NS548;
				when "01010001010" => P_HR_NS <= "0100101" + P_HR_NS549;
				when "01010001011" => P_HR_NS <= "0011101" + P_HR_NS550;
				when "01010001100" => P_HR_NS <= "0100010" + P_HR_NS551;
				when "01010001110" => P_HR_NS <= "0100001" + P_HR_NS552;
				when "01010001111" => P_HR_NS <= "0011111" + P_HR_NS553;
				when "01010010000" => P_HR_NS <= "0100010" + P_HR_NS554;
				when "01010010010" => P_HR_NS <= "0100010" + P_HR_NS555;
				when "01010010011" => P_HR_NS <= "0100100" + P_HR_NS556;
				when "01010010100" => P_HR_NS <= "0100111" + P_HR_NS557;
				when "01010010101" => P_HR_NS <= "0011101" + P_HR_NS558;
				when "01010010111" => P_HR_NS <= "0100000" + P_HR_NS559;
				when "01010011000" => P_HR_NS <= "0011100" + P_HR_NS560;
				when "01010011001" => P_HR_NS <= "0100001" + P_HR_NS561;
				when "01010011011" => P_HR_NS <= "0100100" + P_HR_NS562;
				when "01010011100" => P_HR_NS <= "0100001" + P_HR_NS563;
				when "01010011101" => P_HR_NS <= "0011011" + P_HR_NS564;
				when "01010011111" => P_HR_NS <= "0100010" + P_HR_NS565;
				when "01010100000" => P_HR_NS <= "0011100" + P_HR_NS566;
				when "01010100001" => P_HR_NS <= "0100101" + P_HR_NS567;
				when "01010100011" => P_HR_NS <= "0100110" + P_HR_NS568;
				when "01010100100" => P_HR_NS <= "0100010" + P_HR_NS569;
				when "01010100101" => P_HR_NS <= "0100001" + P_HR_NS570;
				when "01010100111" => P_HR_NS <= "0100000" + P_HR_NS571;
				when "01010101000" => P_HR_NS <= "0011111" + P_HR_NS572;
				when "01010101010" => P_HR_NS <= "0100101" + P_HR_NS573;
				when "01010101011" => P_HR_NS <= "0011100" + P_HR_NS574;
				when "01010101100" => P_HR_NS <= "0011111" + P_HR_NS575;
				when "01010101110" => P_HR_NS <= "0011010" + P_HR_NS576;
				when "01010101111" => P_HR_NS <= "0011100" + P_HR_NS577;
				when "01010110001" => P_HR_NS <= "0011110" + P_HR_NS578;
				when "01010110010" => P_HR_NS <= "0011010" + P_HR_NS579;
				when "01010110011" => P_HR_NS <= "0011010" + P_HR_NS580;
				when "01010110101" => P_HR_NS <= "0100010" + P_HR_NS581;
				when "01010110110" => P_HR_NS <= "0011111" + P_HR_NS582;
				when "01010111000" => P_HR_NS <= "0011111" + P_HR_NS583;
				when "01010111001" => P_HR_NS <= "0011101" + P_HR_NS584;
				when "01010111011" => P_HR_NS <= "0011111" + P_HR_NS585;
				when "01010111100" => P_HR_NS <= "0011011" + P_HR_NS586;
				when "01010111101" => P_HR_NS <= "0011011" + P_HR_NS587;
				when "01010111111" => P_HR_NS <= "0010101" + P_HR_NS588;
				when "01011000000" => P_HR_NS <= "0011001" + P_HR_NS589;
				when "01011000010" => P_HR_NS <= "0011011" + P_HR_NS590;
				when "01011000011" => P_HR_NS <= "0011100" + P_HR_NS591;
				when "01011000101" => P_HR_NS <= "0011111" + P_HR_NS592;
				when "01011000110" => P_HR_NS <= "0010111" + P_HR_NS593;
				when "01011001000" => P_HR_NS <= "0011101" + P_HR_NS594;
				when "01011001001" => P_HR_NS <= "0011010" + P_HR_NS595;
				when "01011001011" => P_HR_NS <= "0011100" + P_HR_NS596;
				when "01011001100" => P_HR_NS <= "0011100" + P_HR_NS597;
				when "01011001110" => P_HR_NS <= "0011010" + P_HR_NS598;
				when "01011001111" => P_HR_NS <= "0010110" + P_HR_NS599;
				when "01011010001" => P_HR_NS <= "0011001" + P_HR_NS600;
				when "01011010011" => P_HR_NS <= "0010111" + P_HR_NS601;
				when "01011010100" => P_HR_NS <= "0010111" + P_HR_NS602;
				when "01011010110" => P_HR_NS <= "0011001" + P_HR_NS603;
				when "01011010111" => P_HR_NS <= "0010101" + P_HR_NS604;
				when "01011011001" => P_HR_NS <= "0010010" + P_HR_NS605;
				when "01011011010" => P_HR_NS <= "0010111" + P_HR_NS606;
				when "01011011100" => P_HR_NS <= "0010011" + P_HR_NS607;
				when "01011011110" => P_HR_NS <= "0010101" + P_HR_NS608;
				when "01011011111" => P_HR_NS <= "0010101" + P_HR_NS609;
				when "01011100001" => P_HR_NS <= "0010110" + P_HR_NS610;
				when "01011100010" => P_HR_NS <= "0010101" + P_HR_NS611;
				when "01011100100" => P_HR_NS <= "0010100" + P_HR_NS612;
				when "01011100110" => P_HR_NS <= "0010011" + P_HR_NS613;
				when "01011100111" => P_HR_NS <= "0001110" + P_HR_NS614;
				when "01011101001" => P_HR_NS <= "0010011" + P_HR_NS615;
				when "01011101011" => P_HR_NS <= "0010001" + P_HR_NS616;
				when "01011101100" => P_HR_NS <= "0001111" + P_HR_NS617;
				when "01011101110" => P_HR_NS <= "0001111" + P_HR_NS618;
				when "01011110000" => P_HR_NS <= "0001011" + P_HR_NS619;
				when "01011110001" => P_HR_NS <= "0010011" + P_HR_NS620;
				when "01011110011" => P_HR_NS <= "0001101" + P_HR_NS621;
				when "01011110101" => P_HR_NS <= "0001100" + P_HR_NS622;
				when "01011110110" => P_HR_NS <= "0010001" + P_HR_NS623;
				when "01011111000" => P_HR_NS <= "0000110" + P_HR_NS624;
				when "01011111010" => P_HR_NS <= "0001100" + P_HR_NS625;
				when "01011111100" => P_HR_NS <= "0001101" + P_HR_NS626;
				when "01011111101" => P_HR_NS <= "0001111" + P_HR_NS627;
				when "01011111111" => P_HR_NS <= "0001011" + P_HR_NS628;
				when "01100000001" => P_HR_NS <= "0001101" + P_HR_NS629;
				when "01100000011" => P_HR_NS <= "0001011" + P_HR_NS630;
				when "01100000100" => P_HR_NS <= "0001101" + P_HR_NS631;
				when "01100000110" => P_HR_NS <= "0001111" + P_HR_NS632;
				when "01100001000" => P_HR_NS <= "0001010" + P_HR_NS633;
				when "01100001010" => P_HR_NS <= "0001011" + P_HR_NS634;
				when "01100001100" => P_HR_NS <= "0001101" + P_HR_NS635;
				when "01100001101" => P_HR_NS <= "0001001" + P_HR_NS636;
				when "01100001111" => P_HR_NS <= "0000110" + P_HR_NS637;
				when "01100010001" => P_HR_NS <= "0001111" + P_HR_NS638;
				when "01100010011" => P_HR_NS <= "0001110" + P_HR_NS639;
				when "01100010101" => P_HR_NS <= "0001001" + P_HR_NS640;
				when "01100010111" => P_HR_NS <= "0001011" + P_HR_NS641;
				when "01100011000" => P_HR_NS <= "0001001" + P_HR_NS642;
				when "01100011010" => P_HR_NS <= "0001000" + P_HR_NS643;
				when "01100011100" => P_HR_NS <= "0001001" + P_HR_NS644;
				when "01100011110" => P_HR_NS <= "0001000" + P_HR_NS645;
				when "01100100000" => P_HR_NS <= "0000111" + P_HR_NS646;
				when "01100100010" => P_HR_NS <= "0000110" + P_HR_NS647;
				when "01100100100" => P_HR_NS <= "0001001" + P_HR_NS648;
				when "01100100110" => P_HR_NS <= "0001000" + P_HR_NS649;
				when "01100101000" => P_HR_NS <= "0000111" + P_HR_NS650;
				when "01100101010" => P_HR_NS <= "0000111" + P_HR_NS651;
				when "01100101100" => P_HR_NS <= "0001000" + P_HR_NS652;
				when "01100101110" => P_HR_NS <= "0000110" + P_HR_NS653;
				when "01100110000" => P_HR_NS <= "0000100" + P_HR_NS654;
				when "01100110010" => P_HR_NS <= "0001000" + P_HR_NS655;
				when "01100110100" => P_HR_NS <= "0000101" + P_HR_NS656;
				when "01100110110" => P_HR_NS <= "0000111" + P_HR_NS657;
				when "01100111000" => P_HR_NS <= "0000110" + P_HR_NS658;
				when "01100111010" => P_HR_NS <= "0000111" + P_HR_NS659;
				when "01100111100" => P_HR_NS <= "0000101" + P_HR_NS660;
				when "01100111110" => P_HR_NS <= "0001010" + P_HR_NS661;
				when "01101000000" => P_HR_NS <= "0000101" + P_HR_NS662;
				when "01101000010" => P_HR_NS <= "0000101" + P_HR_NS663;
				when "01101000100" => P_HR_NS <= "0000101" + P_HR_NS664;
				when "01101000110" => P_HR_NS <= "0000011" + P_HR_NS665;
				when "01101001000" => P_HR_NS <= "0000011" + P_HR_NS666;
				when "01101001010" => P_HR_NS <= "0000100" + P_HR_NS667;
				when "01101001100" => P_HR_NS <= "0000110" + P_HR_NS668;
				when "01101001110" => P_HR_NS <= "0000110" + P_HR_NS669;
				when "01101010000" => P_HR_NS <= "0000110" + P_HR_NS670;
				when "01101010011" => P_HR_NS <= "0000011" + P_HR_NS671;
				when "01101010101" => P_HR_NS <= "0000100" + P_HR_NS672;
				when "01101010111" => P_HR_NS <= "0000100" + P_HR_NS673;
				when "01101011001" => P_HR_NS <= "0000101" + P_HR_NS674;
				when "01101011011" => P_HR_NS <= "0000011" + P_HR_NS675;
				when "01101011110" => P_HR_NS <= "0000110" + P_HR_NS676;
				when "01101100000" => P_HR_NS <= "0000011" + P_HR_NS677;
				when "01101100010" => P_HR_NS <= "0000101" + P_HR_NS678;
				when "01101100100" => P_HR_NS <= "0000011" + P_HR_NS679;
				when "01101100110" => P_HR_NS <= "0000010" + P_HR_NS680;
				when "01101101001" => P_HR_NS <= "0000011" + P_HR_NS681;
				when "01101101011" => P_HR_NS <= "0000011" + P_HR_NS682;
				when "01101101101" => P_HR_NS <= "0000010" + P_HR_NS683;
				when "01101110000" => P_HR_NS <= "0000011" + P_HR_NS684;
				when "01101110010" => P_HR_NS <= "0000011" + P_HR_NS685;
				when "01101110100" => P_HR_NS <= "0000100" + P_HR_NS686;
				when "01101110111" => P_HR_NS <= "0000011" + P_HR_NS687;
				when "01101111001" => P_HR_NS <= "0000011" + P_HR_NS688;
				when "01101111011" => P_HR_NS <= "0000001" + P_HR_NS689;
				when "01101111110" => P_HR_NS <= "0000001" + P_HR_NS690;
				when "01110000000" => P_HR_NS <= "0000001" + P_HR_NS691;
				when "01110000010" => P_HR_NS <= "0000001" + P_HR_NS692;
				when "01110000101" => P_HR_NS <= "0000010" + P_HR_NS693;
				when "01110000111" => P_HR_NS <= "0000010" + P_HR_NS694;
				when "01110001010" => P_HR_NS <= "0000010" + P_HR_NS695;
				when "01110001100" => P_HR_NS <= "0000010" + P_HR_NS696;
				when "01110001111" => P_HR_NS <= "0000010" + P_HR_NS697;
				when "01110010001" => P_HR_NS <= "0000010" + P_HR_NS698;
				when "01110010100" => P_HR_NS <= "0000010" + P_HR_NS699;
				when "01110010110" => P_HR_NS <= "0000010" + P_HR_NS700;
				when "01110011001" => P_HR_NS <= "0000010" + P_HR_NS701;
				when "01110011011" => P_HR_NS <= "0000001" + P_HR_NS702;
				when "01110011110" => P_HR_NS <= "0000010" + P_HR_NS703;
				when "01110100000" => P_HR_NS <= "0000001" + P_HR_NS704;
				when "01110100011" => P_HR_NS <= "0000010" + P_HR_NS705;
				when "01110101000" => P_HR_NS <= "0000001" + P_HR_NS706;
				when "01110101011" => P_HR_NS <= "0000001" + P_HR_NS707;
				when "01110101101" => P_HR_NS <= "0000001" + P_HR_NS708;
				when "01110110000" => P_HR_NS <= "0000001" + P_HR_NS709;
				when "01110110101" => P_HR_NS <= "0000001" + P_HR_NS710;
				when "01110111000" => P_HR_NS <= "0000001" + P_HR_NS711;
				when "01110111011" => P_HR_NS <= "0000001" + P_HR_NS712;
				when "01110111101" => P_HR_NS <= "0000001" + P_HR_NS713;
				when "01111001011" => P_HR_NS <= "0000001" + P_HR_NS714;
				when "01111010001" => P_HR_NS <= "0000001" + P_HR_NS715;
				when "01111011001" => P_HR_NS <= "0000001" + P_HR_NS716;
				when "01111011100" => P_HR_NS <= "0000001" + P_HR_NS717;
				when "01111100101" => P_HR_NS <= "0000001" + P_HR_NS718;
				when "10010000011" => P_HR_NS <= "0000001" + P_HR_NS719;
				when "10010011011" => P_HR_NS <= "0000001" + P_HR_NS720;
				when "10100101011" => P_HR_NS <= "0000001" + P_HR_NS721;
				when "10101100001" => P_HR_NS <= "0000001" + P_HR_NS722;
				when "10101100111" => P_HR_NS <= "0000001" + P_HR_NS723;
				when "10110011100" => P_HR_NS <= "0000001" + P_HR_NS724;
				when "11100000101" => P_HR_NS <= "0000001" + P_HR_NS725;
				when "11110101101" => P_HR_NS <= "0000001" + P_HR_NS726;
				when others            => P_HR_NS <= "000000000001";
			end case;

			case eda is
				when "00000010" => P_EDA_NS <= "000000001" + P_EDA_NS1;
				when "00000011" => P_EDA_NS <= "000000001" + P_EDA_NS2;
				when "00000100" => P_EDA_NS <= "000110111" + P_EDA_NS3;
				when "00000101" => P_EDA_NS <= "001000010" + P_EDA_NS4;
				when "00000110" => P_EDA_NS <= "101010110" + P_EDA_NS5;
				when "00000111" => P_EDA_NS <= "100000111" + P_EDA_NS6;
				when "00001000" => P_EDA_NS <= "111000001" + P_EDA_NS7;
				when "00001001" => P_EDA_NS <= "000111010" + P_EDA_NS8;
				when "00001010" => P_EDA_NS <= "100110100" + P_EDA_NS9;
				when "00001011" => P_EDA_NS <= "011101100" + P_EDA_NS10;
				when "00001100" => P_EDA_NS <= "010101100" + P_EDA_NS11;
				when "00001101" => P_EDA_NS <= "100010011" + P_EDA_NS12;
				when "00001110" => P_EDA_NS <= "011110100" + P_EDA_NS13;
				when "00001111" => P_EDA_NS <= "011011100" + P_EDA_NS14;
				when "00010000" => P_EDA_NS <= "010100111" + P_EDA_NS15;
				when "00010001" => P_EDA_NS <= "010100101" + P_EDA_NS16;
				when "00010010" => P_EDA_NS <= "000101110" + P_EDA_NS17;
				when "00010011" => P_EDA_NS <= "101011111" + P_EDA_NS18;
				when "00010100" => P_EDA_NS <= "010100111" + P_EDA_NS19;
				when "00010101" => P_EDA_NS <= "001110010" + P_EDA_NS20;
				when "00010110" => P_EDA_NS <= "011111101" + P_EDA_NS21;
				when "00010111" => P_EDA_NS <= "111011000" + P_EDA_NS22;
				when "00011000" => P_EDA_NS <= "101111101" + P_EDA_NS23;
				when "00011001" => P_EDA_NS <= "001010011" + P_EDA_NS24;
				when "00011010" => P_EDA_NS <= "000101010" + P_EDA_NS25;
				when "00011011" => P_EDA_NS <= "000001111" + P_EDA_NS26;
				when "00011100" => P_EDA_NS <= "010110000" + P_EDA_NS27;
				when "00011101" => P_EDA_NS <= "010001011" + P_EDA_NS28;
				when "00011110" => P_EDA_NS <= "111110001" + P_EDA_NS29;
				when "00011111" => P_EDA_NS <= "011010000" + P_EDA_NS30;
				when "00100000" => P_EDA_NS <= "010011001" + P_EDA_NS31;
				when "00100001" => P_EDA_NS <= "000101001" + P_EDA_NS32;
				when "00100010" => P_EDA_NS <= "000001110" + P_EDA_NS33;
				when "00100011" => P_EDA_NS <= "000001100" + P_EDA_NS34;
				when "00100100" => P_EDA_NS <= "000001101" + P_EDA_NS35;
				when "00100101" => P_EDA_NS <= "000001100" + P_EDA_NS36;
				when "00100110" => P_EDA_NS <= "000001010" + P_EDA_NS37;
				when "00100111" => P_EDA_NS <= "000000111" + P_EDA_NS38;
				when "00101000" => P_EDA_NS <= "000001100" + P_EDA_NS39;
				when "00101001" => P_EDA_NS <= "000010100" + P_EDA_NS40;
				when "00101010" => P_EDA_NS <= "001001000" + P_EDA_NS41;
				when "00101011" => P_EDA_NS <= "010010001" + P_EDA_NS42;
				when "00101100" => P_EDA_NS <= "010011000" + P_EDA_NS43;
				when "00101101" => P_EDA_NS <= "000110110" + P_EDA_NS44;
				when "00101110" => P_EDA_NS <= "000110110" + P_EDA_NS45;
				when "00101111" => P_EDA_NS <= "000101110" + P_EDA_NS46;
				when "00110000" => P_EDA_NS <= "011110101" + P_EDA_NS47;
				when "00110001" => P_EDA_NS <= "011001010" + P_EDA_NS48;
				when "00110010" => P_EDA_NS <= "100001010" + P_EDA_NS49;
				when "00110011" => P_EDA_NS <= "011100101" + P_EDA_NS50;
				when "00110100" => P_EDA_NS <= "011010110" + P_EDA_NS51;
				when "00110101" => P_EDA_NS <= "010001000" + P_EDA_NS52;
				when "00110110" => P_EDA_NS <= "000111111" + P_EDA_NS53;
				when "00110111" => P_EDA_NS <= "000100011" + P_EDA_NS54;
				when "00111000" => P_EDA_NS <= "001000001" + P_EDA_NS55;
				when "00111001" => P_EDA_NS <= "011010100" + P_EDA_NS56;
				when "00111010" => P_EDA_NS <= "001011001" + P_EDA_NS57;
				when "00111011" => P_EDA_NS <= "000111000" + P_EDA_NS58;
				when "00111100" => P_EDA_NS <= "001000101" + P_EDA_NS59;
				when "00111101" => P_EDA_NS <= "001010110" + P_EDA_NS60;
				when "00111110" => P_EDA_NS <= "000110010" + P_EDA_NS61;
				when "00111111" => P_EDA_NS <= "000111001" + P_EDA_NS62;
				when "01000000" => P_EDA_NS <= "000101001" + P_EDA_NS63;
				when "01000001" => P_EDA_NS <= "000101100" + P_EDA_NS64;
				when "01000010" => P_EDA_NS <= "001001101" + P_EDA_NS65;
				when "01000011" => P_EDA_NS <= "000110011" + P_EDA_NS66;
				when "01000100" => P_EDA_NS <= "000011111" + P_EDA_NS67;
				when "01000101" => P_EDA_NS <= "000011011" + P_EDA_NS68;
				when "01000110" => P_EDA_NS <= "000100010" + P_EDA_NS69;
				when "01000111" => P_EDA_NS <= "000010001" + P_EDA_NS70;
				when "01001000" => P_EDA_NS <= "000001011" + P_EDA_NS71;
				when "01001001" => P_EDA_NS <= "000001010" + P_EDA_NS72;
				when "01001010" => P_EDA_NS <= "000001001" + P_EDA_NS73;
				when "01001011" => P_EDA_NS <= "000001001" + P_EDA_NS74;
				when "01001100" => P_EDA_NS <= "000001011" + P_EDA_NS75;
				when "01001101" => P_EDA_NS <= "000001000" + P_EDA_NS76;
				when "01001110" => P_EDA_NS <= "000000110" + P_EDA_NS77;
				when "01001111" => P_EDA_NS <= "000001101" + P_EDA_NS78;
				when "01010000" => P_EDA_NS <= "000001001" + P_EDA_NS79;
				when "01010001" => P_EDA_NS <= "000000010" + P_EDA_NS80;
				when "01010010" => P_EDA_NS <= "000000100" + P_EDA_NS81;
				when "01010011" => P_EDA_NS <= "000000011" + P_EDA_NS82;
				when "01010100" => P_EDA_NS <= "000000010" + P_EDA_NS83;
				when "01010101" => P_EDA_NS <= "000000010" + P_EDA_NS84;
				when "01010110" => P_EDA_NS <= "000000010" + P_EDA_NS85;
				when "01010111" => P_EDA_NS <= "000000010" + P_EDA_NS86;
				when "01011000" => P_EDA_NS <= "000000001" + P_EDA_NS87;
				when "01011001" => P_EDA_NS <= "001010101" + P_EDA_NS88;
				when "01011010" => P_EDA_NS <= "001100110" + P_EDA_NS89;
				when "01011011" => P_EDA_NS <= "000100100" + P_EDA_NS90;
				when "01011100" => P_EDA_NS <= "001100011" + P_EDA_NS91;
				when "01011101" => P_EDA_NS <= "001000010" + P_EDA_NS92;
				when "01011110" => P_EDA_NS <= "001000000" + P_EDA_NS93;
				when "01011111" => P_EDA_NS <= "000110110" + P_EDA_NS94;
				when "01100000" => P_EDA_NS <= "000011110" + P_EDA_NS95;
				when "01100001" => P_EDA_NS <= "000001011" + P_EDA_NS96;
				when "01100010" => P_EDA_NS <= "000001110" + P_EDA_NS97;
				when "01100011" => P_EDA_NS <= "000011101" + P_EDA_NS98;
				when "01100100" => P_EDA_NS <= "000001110" + P_EDA_NS99;
				when "01100101" => P_EDA_NS <= "000010001" + P_EDA_NS100;
				when "01100110" => P_EDA_NS <= "000001110" + P_EDA_NS101;
				when "01100111" => P_EDA_NS <= "000001110" + P_EDA_NS102;
				when "01101000" => P_EDA_NS <= "000010101" + P_EDA_NS103;
				when "01101001" => P_EDA_NS <= "000001001" + P_EDA_NS104;
				when "01101010" => P_EDA_NS <= "000000111" + P_EDA_NS105;
				when "01101011" => P_EDA_NS <= "000001010" + P_EDA_NS106;
				when "01101100" => P_EDA_NS <= "000000001" + P_EDA_NS107;
				when "10101110" => P_EDA_NS <= "000000010" + P_EDA_NS108;
				when "10101111" => P_EDA_NS <= "000000111" + P_EDA_NS109;
				when "10110000" => P_EDA_NS <= "000000100" + P_EDA_NS110;
				when others    => P_EDA_NS <= "000000000001";
			end case;
			not_stress_score <= P_TEMP_NS * P_NOT_STRESS * P_EDA_NS * P_HR_NS;
			
			--not_stress_score <= P_TEMP_NS * P_NOT_STRESS * P_EDA_NS * P_HR_NS;
		elsif (state = TRAINING_NS) then
			
			case temp is
				when "011100000" => P_TEMP_NS1 <= P_TEMP_NS1 + T_N_STRESS;
				when "011100001" => P_TEMP_NS2 <= P_TEMP_NS2 + T_N_STRESS;
				when "011100010" => P_TEMP_NS3 <= P_TEMP_NS3 + T_N_STRESS;
				when "011100011" => P_TEMP_NS4 <= P_TEMP_NS4 + T_N_STRESS;
				when "011100100" => P_TEMP_NS5 <= P_TEMP_NS5 + T_N_STRESS;
				when "011100101" => P_TEMP_NS6 <= P_TEMP_NS6 + T_N_STRESS;
				when "011100110" => P_TEMP_NS7 <= P_TEMP_NS7 + T_N_STRESS;
				when "011100111" => P_TEMP_NS8 <= P_TEMP_NS8 + T_N_STRESS;
				when "011101000" => P_TEMP_NS9 <= P_TEMP_NS9 + T_N_STRESS;
				when "011101001" => P_TEMP_NS10 <= P_TEMP_NS10 + T_N_STRESS;
				when "011101010" => P_TEMP_NS11 <= P_TEMP_NS11 + T_N_STRESS;
				when "011101011" => P_TEMP_NS12 <= P_TEMP_NS12 + T_N_STRESS;
				when "011101100" => P_TEMP_NS13 <= P_TEMP_NS13 + T_N_STRESS;
				when "011101101" => P_TEMP_NS14 <= P_TEMP_NS14 + T_N_STRESS;
				when "011101110" => P_TEMP_NS15 <= P_TEMP_NS15 + T_N_STRESS;
				when "011101111" => P_TEMP_NS16 <= P_TEMP_NS16 + T_N_STRESS;
				when "011110000" => P_TEMP_NS17 <= P_TEMP_NS17 + T_N_STRESS;
				when "011110001" => P_TEMP_NS18 <= P_TEMP_NS18 + T_N_STRESS;
				when "011110010" => P_TEMP_NS19 <= P_TEMP_NS19 + T_N_STRESS;
				when "011110011" => P_TEMP_NS20 <= P_TEMP_NS20 + T_N_STRESS;
				when "011110100" => P_TEMP_NS21 <= P_TEMP_NS21 + T_N_STRESS;
				when "011110101" => P_TEMP_NS22 <= P_TEMP_NS22 + T_N_STRESS;
				when "011110110" => P_TEMP_NS23 <= P_TEMP_NS23 + T_N_STRESS;
				when "011110111" => P_TEMP_NS24 <= P_TEMP_NS24 + T_N_STRESS;
				when "011111000" => P_TEMP_NS25 <= P_TEMP_NS25 + T_N_STRESS;
				when "011111001" => P_TEMP_NS26 <= P_TEMP_NS26 + T_N_STRESS;
				when "011111010" => P_TEMP_NS27 <= P_TEMP_NS27 + T_N_STRESS;
				when "011111011" => P_TEMP_NS28 <= P_TEMP_NS28 + T_N_STRESS;
				when "011111100" => P_TEMP_NS29 <= P_TEMP_NS29 + T_N_STRESS;
				when "011111101" => P_TEMP_NS30 <= P_TEMP_NS30 + T_N_STRESS;
				when "011111110" => P_TEMP_NS31 <= P_TEMP_NS31 + T_N_STRESS;
				when "011111111" => P_TEMP_NS32 <= P_TEMP_NS32 + T_N_STRESS;
				when "100000000" => P_TEMP_NS33 <= P_TEMP_NS33 + T_N_STRESS;
				when "100000001" => P_TEMP_NS34 <= P_TEMP_NS34 + T_N_STRESS;
				when "100000010" => P_TEMP_NS35 <= P_TEMP_NS35 + T_N_STRESS;
				when "100000011" => P_TEMP_NS36 <= P_TEMP_NS36 + T_N_STRESS;
				when "100000100" => P_TEMP_NS37 <= P_TEMP_NS37 + T_N_STRESS;
				when "100000101" => P_TEMP_NS38 <= P_TEMP_NS38 + T_N_STRESS;
				when "100000110" => P_TEMP_NS39 <= P_TEMP_NS39 + T_N_STRESS;
				when "100000111" => P_TEMP_NS40 <= P_TEMP_NS40 + T_N_STRESS;
				when "100001000" => P_TEMP_NS41 <= P_TEMP_NS41 + T_N_STRESS;
				when "100001001" => P_TEMP_NS42 <= P_TEMP_NS42 + T_N_STRESS;
				when "100001010" => P_TEMP_NS43 <= P_TEMP_NS43 + T_N_STRESS;
				when "100001011" => P_TEMP_NS44 <= P_TEMP_NS44 + T_N_STRESS;
				when "100001100" => P_TEMP_NS45 <= P_TEMP_NS45 + T_N_STRESS;
				when "100001101" => P_TEMP_NS46 <= P_TEMP_NS46 + T_N_STRESS;
				when "100001110" => P_TEMP_NS47 <= P_TEMP_NS47 + T_N_STRESS;
				when "100001111" => P_TEMP_NS48 <= P_TEMP_NS48 + T_N_STRESS;
				when "100010000" => P_TEMP_NS49 <= P_TEMP_NS49 + T_N_STRESS;
				when "100010001" => P_TEMP_NS50 <= P_TEMP_NS50 + T_N_STRESS;
				when "100010010" => P_TEMP_NS51 <= P_TEMP_NS51 + T_N_STRESS;
				when "100010011" => P_TEMP_NS52 <= P_TEMP_NS52 + T_N_STRESS;
				when "100010100" => P_TEMP_NS53 <= P_TEMP_NS53 + T_N_STRESS;
				when "100010101" => P_TEMP_NS54 <= P_TEMP_NS54 + T_N_STRESS;
				when "100010110" => P_TEMP_NS55 <= P_TEMP_NS55 + T_N_STRESS;
				when "100010111" => P_TEMP_NS56 <= P_TEMP_NS56 + T_N_STRESS;
				when "100011000" => P_TEMP_NS57 <= P_TEMP_NS57 + T_N_STRESS;
				when "100011001" => P_TEMP_NS58 <= P_TEMP_NS58 + T_N_STRESS;
				when "100011010" => P_TEMP_NS59 <= P_TEMP_NS59 + T_N_STRESS;
				when "100011011" => P_TEMP_NS60 <= P_TEMP_NS60 + T_N_STRESS;
				when "100011100" => P_TEMP_NS61 <= P_TEMP_NS61 + T_N_STRESS;
				when "100011101" => P_TEMP_NS62 <= P_TEMP_NS62 + T_N_STRESS;
				when "100011110" => P_TEMP_NS63 <= P_TEMP_NS63 + T_N_STRESS;
				when  others     => null;
			end case;	

			case hr is
                when "00000000001" => P_HR_NS1 <= P_HR_NS1 + T_N_STRESS;
                when "00000000011" => P_HR_NS2 <= P_HR_NS2 + T_N_STRESS;
                when "00000000100" => P_HR_NS3 <= P_HR_NS3 + T_N_STRESS;
                when "00000000111" => P_HR_NS4 <= P_HR_NS4 + T_N_STRESS;
                when "00000001000" => P_HR_NS5 <= P_HR_NS5 + T_N_STRESS;
                when "00000001001" => P_HR_NS6 <= P_HR_NS6 + T_N_STRESS;
                when "00000001010" => P_HR_NS7 <= P_HR_NS7 + T_N_STRESS;
                when "00000001100" => P_HR_NS8 <= P_HR_NS8 + T_N_STRESS;
                when "00000001101" => P_HR_NS9 <= P_HR_NS9 + T_N_STRESS;
                when "00000001110" => P_HR_NS10 <= P_HR_NS10 + T_N_STRESS;
                when "00000001111" => P_HR_NS11 <= P_HR_NS11 + T_N_STRESS;
                when "00000010000" => P_HR_NS12 <= P_HR_NS12 + T_N_STRESS;
                when "00000010001" => P_HR_NS13 <= P_HR_NS13 + T_N_STRESS;
                when "00000010010" => P_HR_NS14 <= P_HR_NS14 + T_N_STRESS;
                when "00000010011" => P_HR_NS15 <= P_HR_NS15 + T_N_STRESS;
                when "00000010101" => P_HR_NS16 <= P_HR_NS16 + T_N_STRESS;
                when "00000010110" => P_HR_NS17 <= P_HR_NS17 + T_N_STRESS;
                when "00000011100" => P_HR_NS18 <= P_HR_NS18 + T_N_STRESS;
                when "00000011101" => P_HR_NS19 <= P_HR_NS19 + T_N_STRESS;
                when "00000011110" => P_HR_NS20 <= P_HR_NS20 + T_N_STRESS;
                when "00000011111" => P_HR_NS21 <= P_HR_NS21 + T_N_STRESS;
                when "00000100000" => P_HR_NS22 <= P_HR_NS22 + T_N_STRESS;
                when "00000100010" => P_HR_NS23 <= P_HR_NS23 + T_N_STRESS;
                when "00000100110" => P_HR_NS24 <= P_HR_NS24 + T_N_STRESS;
                when "00000100111" => P_HR_NS25 <= P_HR_NS25 + T_N_STRESS;
                when "00000101000" => P_HR_NS26 <= P_HR_NS26 + T_N_STRESS;
                when "00000101001" => P_HR_NS27 <= P_HR_NS27 + T_N_STRESS;
                when "00000101010" => P_HR_NS28 <= P_HR_NS28 + T_N_STRESS;
                when "00000101011" => P_HR_NS29 <= P_HR_NS29 + T_N_STRESS;
                when "00000110100" => P_HR_NS30 <= P_HR_NS30 + T_N_STRESS;
                when "00000110101" => P_HR_NS31 <= P_HR_NS31 + T_N_STRESS;
                when "00000111000" => P_HR_NS32 <= P_HR_NS32 + T_N_STRESS;
                when "00000111010" => P_HR_NS33 <= P_HR_NS33 + T_N_STRESS;
                when "00000111100" => P_HR_NS34 <= P_HR_NS34 + T_N_STRESS;
                when "00001000001" => P_HR_NS35 <= P_HR_NS35 + T_N_STRESS;
                when "00001000011" => P_HR_NS36 <= P_HR_NS36 + T_N_STRESS;
                when "00001000100" => P_HR_NS37 <= P_HR_NS37 + T_N_STRESS;
                when "00001000110" => P_HR_NS38 <= P_HR_NS38 + T_N_STRESS;
                when "00001001000" => P_HR_NS39 <= P_HR_NS39 + T_N_STRESS;
                when "00001001100" => P_HR_NS40 <= P_HR_NS40 + T_N_STRESS;
                when "00001001101" => P_HR_NS41 <= P_HR_NS41 + T_N_STRESS;
                when "00001001110" => P_HR_NS42 <= P_HR_NS42 + T_N_STRESS;
                when "00001001111" => P_HR_NS43 <= P_HR_NS43 + T_N_STRESS;
                when "00001010011" => P_HR_NS44 <= P_HR_NS44 + T_N_STRESS;
                when "00001010101" => P_HR_NS45 <= P_HR_NS45 + T_N_STRESS;
                when "00001010110" => P_HR_NS46 <= P_HR_NS46 + T_N_STRESS;
                when "00001011000" => P_HR_NS47 <= P_HR_NS47 + T_N_STRESS;
                when "00001011001" => P_HR_NS48 <= P_HR_NS48 + T_N_STRESS;
                when "00001011010" => P_HR_NS49 <= P_HR_NS49 + T_N_STRESS;
                when "00001011100" => P_HR_NS50 <= P_HR_NS50 + T_N_STRESS;
                when "00001011111" => P_HR_NS51 <= P_HR_NS51 + T_N_STRESS;
                when "00001100000" => P_HR_NS52 <= P_HR_NS52 + T_N_STRESS;
                when "00001100001" => P_HR_NS53 <= P_HR_NS53 + T_N_STRESS;
                when "00001100101" => P_HR_NS54 <= P_HR_NS54 + T_N_STRESS;
                when "00001101000" => P_HR_NS55 <= P_HR_NS55 + T_N_STRESS;
                when "00001101001" => P_HR_NS56 <= P_HR_NS56 + T_N_STRESS;
                when "00001101011" => P_HR_NS57 <= P_HR_NS57 + T_N_STRESS;
                when "00001101100" => P_HR_NS58 <= P_HR_NS58 + T_N_STRESS;
                when "00001101110" => P_HR_NS59 <= P_HR_NS59 + T_N_STRESS;
                when "00001101111" => P_HR_NS60 <= P_HR_NS60 + T_N_STRESS;
                when "00001110000" => P_HR_NS61 <= P_HR_NS61 + T_N_STRESS;
                when "00001110001" => P_HR_NS62 <= P_HR_NS62 + T_N_STRESS;
                when "00001110010" => P_HR_NS63 <= P_HR_NS63 + T_N_STRESS;
                when "00001110101" => P_HR_NS64 <= P_HR_NS64 + T_N_STRESS;
                when "00001110110" => P_HR_NS65 <= P_HR_NS65 + T_N_STRESS;
                when "00001111000" => P_HR_NS66 <= P_HR_NS66 + T_N_STRESS;
                when "00001111011" => P_HR_NS67 <= P_HR_NS67 + T_N_STRESS;
                when "00001111110" => P_HR_NS68 <= P_HR_NS68 + T_N_STRESS;
                when "00001111111" => P_HR_NS69 <= P_HR_NS69 + T_N_STRESS;
                when "00010000000" => P_HR_NS70 <= P_HR_NS70 + T_N_STRESS;
                when "00010000010" => P_HR_NS71 <= P_HR_NS71 + T_N_STRESS;
                when "00010000100" => P_HR_NS72 <= P_HR_NS72 + T_N_STRESS;
                when "00010000101" => P_HR_NS73 <= P_HR_NS73 + T_N_STRESS;
                when "00010000110" => P_HR_NS74 <= P_HR_NS74 + T_N_STRESS;
                when "00010000111" => P_HR_NS75 <= P_HR_NS75 + T_N_STRESS;
                when "00010001001" => P_HR_NS76 <= P_HR_NS76 + T_N_STRESS;
                when "00010001010" => P_HR_NS77 <= P_HR_NS77 + T_N_STRESS;
                when "00010001011" => P_HR_NS78 <= P_HR_NS78 + T_N_STRESS;
                when "00010001100" => P_HR_NS79 <= P_HR_NS79 + T_N_STRESS;
                when "00010001101" => P_HR_NS80 <= P_HR_NS80 + T_N_STRESS;
                when "00010001111" => P_HR_NS81 <= P_HR_NS81 + T_N_STRESS;
                when "00010010000" => P_HR_NS82 <= P_HR_NS82 + T_N_STRESS;
                when "00010010001" => P_HR_NS83 <= P_HR_NS83 + T_N_STRESS;
                when "00010010010" => P_HR_NS84 <= P_HR_NS84 + T_N_STRESS;
                when "00010010011" => P_HR_NS85 <= P_HR_NS85 + T_N_STRESS;
                when "00010010100" => P_HR_NS86 <= P_HR_NS86 + T_N_STRESS;
                when "00010010101" => P_HR_NS87 <= P_HR_NS87 + T_N_STRESS;
                when "00010010110" => P_HR_NS88 <= P_HR_NS88 + T_N_STRESS;
                when "00010010111" => P_HR_NS89 <= P_HR_NS89 + T_N_STRESS;
                when "00010011001" => P_HR_NS90 <= P_HR_NS90 + T_N_STRESS;
                when "00010011100" => P_HR_NS91 <= P_HR_NS91 + T_N_STRESS;
                when "00010011110" => P_HR_NS92 <= P_HR_NS92 + T_N_STRESS;
                when "00010011111" => P_HR_NS93 <= P_HR_NS93 + T_N_STRESS;
                when "00010100001" => P_HR_NS94 <= P_HR_NS94 + T_N_STRESS;
                when "00010100010" => P_HR_NS95 <= P_HR_NS95 + T_N_STRESS;
                when "00010100011" => P_HR_NS96 <= P_HR_NS96 + T_N_STRESS;
                when "00010100100" => P_HR_NS97 <= P_HR_NS97 + T_N_STRESS;
                when "00010100101" => P_HR_NS98 <= P_HR_NS98 + T_N_STRESS;
                when "00010100110" => P_HR_NS99 <= P_HR_NS99 + T_N_STRESS;
                when "00010100111" => P_HR_NS100 <= P_HR_NS100 + T_N_STRESS;
                when "00010101000" => P_HR_NS101 <= P_HR_NS101 + T_N_STRESS;
                when "00010101001" => P_HR_NS102 <= P_HR_NS102 + T_N_STRESS;
                when "00010101010" => P_HR_NS103 <= P_HR_NS103 + T_N_STRESS;
                when "00010101011" => P_HR_NS104 <= P_HR_NS104 + T_N_STRESS;
                when "00010101101" => P_HR_NS105 <= P_HR_NS105 + T_N_STRESS;
                when "00010101110" => P_HR_NS106 <= P_HR_NS106 + T_N_STRESS;
                when "00010101111" => P_HR_NS107 <= P_HR_NS107 + T_N_STRESS;
                when "00010110000" => P_HR_NS108 <= P_HR_NS108 + T_N_STRESS;
                when "00010110001" => P_HR_NS109 <= P_HR_NS109 + T_N_STRESS;
                when "00010110010" => P_HR_NS110 <= P_HR_NS110 + T_N_STRESS;
                when "00010110011" => P_HR_NS111 <= P_HR_NS111 + T_N_STRESS;
                when "00010110100" => P_HR_NS112 <= P_HR_NS112 + T_N_STRESS;
                when "00010110101" => P_HR_NS113 <= P_HR_NS113 + T_N_STRESS;
                when "00010110110" => P_HR_NS114 <= P_HR_NS114 + T_N_STRESS;
                when "00010110111" => P_HR_NS115 <= P_HR_NS115 + T_N_STRESS;
                when "00010111000" => P_HR_NS116 <= P_HR_NS116 + T_N_STRESS;
                when "00010111001" => P_HR_NS117 <= P_HR_NS117 + T_N_STRESS;
                when "00010111010" => P_HR_NS118 <= P_HR_NS118 + T_N_STRESS;
                when "00010111011" => P_HR_NS119 <= P_HR_NS119 + T_N_STRESS;
                when "00010111100" => P_HR_NS120 <= P_HR_NS120 + T_N_STRESS;
                when "00010111101" => P_HR_NS121 <= P_HR_NS121 + T_N_STRESS;
                when "00010111110" => P_HR_NS122 <= P_HR_NS122 + T_N_STRESS;
                when "00010111111" => P_HR_NS123 <= P_HR_NS123 + T_N_STRESS;
                when "00011000000" => P_HR_NS124 <= P_HR_NS124 + T_N_STRESS;
                when "00011000001" => P_HR_NS125 <= P_HR_NS125 + T_N_STRESS;
                when "00011000010" => P_HR_NS126 <= P_HR_NS126 + T_N_STRESS;
                when "00011000011" => P_HR_NS127 <= P_HR_NS127 + T_N_STRESS;
                when "00011000100" => P_HR_NS128 <= P_HR_NS128 + T_N_STRESS;
                when "00011000101" => P_HR_NS129 <= P_HR_NS129 + T_N_STRESS;
                when "00011000110" => P_HR_NS130 <= P_HR_NS130 + T_N_STRESS;
                when "00011000111" => P_HR_NS131 <= P_HR_NS131 + T_N_STRESS;
                when "00011001000" => P_HR_NS132 <= P_HR_NS132 + T_N_STRESS;
                when "00011001001" => P_HR_NS133 <= P_HR_NS133 + T_N_STRESS;
                when "00011001010" => P_HR_NS134 <= P_HR_NS134 + T_N_STRESS;
                when "00011001011" => P_HR_NS135 <= P_HR_NS135 + T_N_STRESS;
                when "00011001100" => P_HR_NS136 <= P_HR_NS136 + T_N_STRESS;
                when "00011001101" => P_HR_NS137 <= P_HR_NS137 + T_N_STRESS;
                when "00011001111" => P_HR_NS138 <= P_HR_NS138 + T_N_STRESS;
                when "00011010000" => P_HR_NS139 <= P_HR_NS139 + T_N_STRESS;
                when "00011010001" => P_HR_NS140 <= P_HR_NS140 + T_N_STRESS;
                when "00011010010" => P_HR_NS141 <= P_HR_NS141 + T_N_STRESS;
                when "00011010011" => P_HR_NS142 <= P_HR_NS142 + T_N_STRESS;
                when "00011010100" => P_HR_NS143 <= P_HR_NS143 + T_N_STRESS;
                when "00011010101" => P_HR_NS144 <= P_HR_NS144 + T_N_STRESS;
                when "00011010110" => P_HR_NS145 <= P_HR_NS145 + T_N_STRESS;
                when "00011010111" => P_HR_NS146 <= P_HR_NS146 + T_N_STRESS;
                when "00011011000" => P_HR_NS147 <= P_HR_NS147 + T_N_STRESS;
                when "00011011001" => P_HR_NS148 <= P_HR_NS148 + T_N_STRESS;
                when "00011011011" => P_HR_NS149 <= P_HR_NS149 + T_N_STRESS;
                when "00011100000" => P_HR_NS150 <= P_HR_NS150 + T_N_STRESS;
                when "00011100010" => P_HR_NS151 <= P_HR_NS151 + T_N_STRESS;
                when "00011100011" => P_HR_NS152 <= P_HR_NS152 + T_N_STRESS;
                when "00011100100" => P_HR_NS153 <= P_HR_NS153 + T_N_STRESS;
                when "00011100101" => P_HR_NS154 <= P_HR_NS154 + T_N_STRESS;
                when "00011100110" => P_HR_NS155 <= P_HR_NS155 + T_N_STRESS;
                when "00011100111" => P_HR_NS156 <= P_HR_NS156 + T_N_STRESS;
                when "00011101000" => P_HR_NS157 <= P_HR_NS157 + T_N_STRESS;
                when "00011101001" => P_HR_NS158 <= P_HR_NS158 + T_N_STRESS;
                when "00011101010" => P_HR_NS159 <= P_HR_NS159 + T_N_STRESS;
                when "00011101011" => P_HR_NS160 <= P_HR_NS160 + T_N_STRESS;
                when "00011101101" => P_HR_NS161 <= P_HR_NS161 + T_N_STRESS;
                when "00011101111" => P_HR_NS162 <= P_HR_NS162 + T_N_STRESS;
                when "00011110000" => P_HR_NS163 <= P_HR_NS163 + T_N_STRESS;
                when "00011110011" => P_HR_NS164 <= P_HR_NS164 + T_N_STRESS;
                when "00011110101" => P_HR_NS165 <= P_HR_NS165 + T_N_STRESS;
                when "00011110110" => P_HR_NS166 <= P_HR_NS166 + T_N_STRESS;
                when "00011111000" => P_HR_NS167 <= P_HR_NS167 + T_N_STRESS;
                when "00011111001" => P_HR_NS168 <= P_HR_NS168 + T_N_STRESS;
                when "00011111010" => P_HR_NS169 <= P_HR_NS169 + T_N_STRESS;
                when "00011111011" => P_HR_NS170 <= P_HR_NS170 + T_N_STRESS;
                when "00011111100" => P_HR_NS171 <= P_HR_NS171 + T_N_STRESS;
                when "00011111101" => P_HR_NS172 <= P_HR_NS172 + T_N_STRESS;
                when "00011111110" => P_HR_NS173 <= P_HR_NS173 + T_N_STRESS;
                when "00011111111" => P_HR_NS174 <= P_HR_NS174 + T_N_STRESS;
                when "00100000000" => P_HR_NS175 <= P_HR_NS175 + T_N_STRESS;
                when "00100000001" => P_HR_NS176 <= P_HR_NS176 + T_N_STRESS;
                when "00100000010" => P_HR_NS177 <= P_HR_NS177 + T_N_STRESS;
                when "00100000011" => P_HR_NS178 <= P_HR_NS178 + T_N_STRESS;
                when "00100000100" => P_HR_NS179 <= P_HR_NS179 + T_N_STRESS;
                when "00100000101" => P_HR_NS180 <= P_HR_NS180 + T_N_STRESS;
                when "00100000110" => P_HR_NS181 <= P_HR_NS181 + T_N_STRESS;
                when "00100000111" => P_HR_NS182 <= P_HR_NS182 + T_N_STRESS;
                when "00100001000" => P_HR_NS183 <= P_HR_NS183 + T_N_STRESS;
                when "00100001001" => P_HR_NS184 <= P_HR_NS184 + T_N_STRESS;
                when "00100001010" => P_HR_NS185 <= P_HR_NS185 + T_N_STRESS;
                when "00100001011" => P_HR_NS186 <= P_HR_NS186 + T_N_STRESS;
                when "00100001100" => P_HR_NS187 <= P_HR_NS187 + T_N_STRESS;
                when "00100001101" => P_HR_NS188 <= P_HR_NS188 + T_N_STRESS;
                when "00100001110" => P_HR_NS189 <= P_HR_NS189 + T_N_STRESS;
                when "00100001111" => P_HR_NS190 <= P_HR_NS190 + T_N_STRESS;
                when "00100010000" => P_HR_NS191 <= P_HR_NS191 + T_N_STRESS;
                when "00100010001" => P_HR_NS192 <= P_HR_NS192 + T_N_STRESS;
                when "00100010010" => P_HR_NS193 <= P_HR_NS193 + T_N_STRESS;
                when "00100010011" => P_HR_NS194 <= P_HR_NS194 + T_N_STRESS;
                when "00100010100" => P_HR_NS195 <= P_HR_NS195 + T_N_STRESS;
                when "00100010101" => P_HR_NS196 <= P_HR_NS196 + T_N_STRESS;
                when "00100010110" => P_HR_NS197 <= P_HR_NS197 + T_N_STRESS;
                when "00100010111" => P_HR_NS198 <= P_HR_NS198 + T_N_STRESS;
                when "00100011000" => P_HR_NS199 <= P_HR_NS199 + T_N_STRESS;
                when "00100011001" => P_HR_NS200 <= P_HR_NS200 + T_N_STRESS;
                when "00100011010" => P_HR_NS201 <= P_HR_NS201 + T_N_STRESS;
                when "00100011011" => P_HR_NS202 <= P_HR_NS202 + T_N_STRESS;
                when "00100011100" => P_HR_NS203 <= P_HR_NS203 + T_N_STRESS;
                when "00100011101" => P_HR_NS204 <= P_HR_NS204 + T_N_STRESS;
                when "00100011110" => P_HR_NS205 <= P_HR_NS205 + T_N_STRESS;
                when "00100011111" => P_HR_NS206 <= P_HR_NS206 + T_N_STRESS;
                when "00100100000" => P_HR_NS207 <= P_HR_NS207 + T_N_STRESS;
                when "00100100001" => P_HR_NS208 <= P_HR_NS208 + T_N_STRESS;
                when "00100100010" => P_HR_NS209 <= P_HR_NS209 + T_N_STRESS;
                when "00100100011" => P_HR_NS210 <= P_HR_NS210 + T_N_STRESS;
                when "00100100100" => P_HR_NS211 <= P_HR_NS211 + T_N_STRESS;
                when "00100100101" => P_HR_NS212 <= P_HR_NS212 + T_N_STRESS;
                when "00100100110" => P_HR_NS213 <= P_HR_NS213 + T_N_STRESS;
                when "00100101001" => P_HR_NS214 <= P_HR_NS214 + T_N_STRESS;
                when "00100101010" => P_HR_NS215 <= P_HR_NS215 + T_N_STRESS;
                when "00100101011" => P_HR_NS216 <= P_HR_NS216 + T_N_STRESS;
                when "00100101100" => P_HR_NS217 <= P_HR_NS217 + T_N_STRESS;
                when "00100101101" => P_HR_NS218 <= P_HR_NS218 + T_N_STRESS;
                when "00100101110" => P_HR_NS219 <= P_HR_NS219 + T_N_STRESS;
                when "00100110000" => P_HR_NS220 <= P_HR_NS220 + T_N_STRESS;
                when "00100110010" => P_HR_NS221 <= P_HR_NS221 + T_N_STRESS;
                when "00100110011" => P_HR_NS222 <= P_HR_NS222 + T_N_STRESS;
                when "00100110100" => P_HR_NS223 <= P_HR_NS223 + T_N_STRESS;
                when "00100110110" => P_HR_NS224 <= P_HR_NS224 + T_N_STRESS;
                when "00100111000" => P_HR_NS225 <= P_HR_NS225 + T_N_STRESS;
                when "00100111010" => P_HR_NS226 <= P_HR_NS226 + T_N_STRESS;
                when "00100111011" => P_HR_NS227 <= P_HR_NS227 + T_N_STRESS;
                when "00100111100" => P_HR_NS228 <= P_HR_NS228 + T_N_STRESS;
                when "00100111110" => P_HR_NS229 <= P_HR_NS229 + T_N_STRESS;
                when "00100111111" => P_HR_NS230 <= P_HR_NS230 + T_N_STRESS;
                when "00101000000" => P_HR_NS231 <= P_HR_NS231 + T_N_STRESS;
                when "00101000010" => P_HR_NS232 <= P_HR_NS232 + T_N_STRESS;
                when "00101000011" => P_HR_NS233 <= P_HR_NS233 + T_N_STRESS;
                when "00101000100" => P_HR_NS234 <= P_HR_NS234 + T_N_STRESS;
                when "00101000101" => P_HR_NS235 <= P_HR_NS235 + T_N_STRESS;
                when "00101000110" => P_HR_NS236 <= P_HR_NS236 + T_N_STRESS;
                when "00101000111" => P_HR_NS237 <= P_HR_NS237 + T_N_STRESS;
                when "00101001000" => P_HR_NS238 <= P_HR_NS238 + T_N_STRESS;
                when "00101001011" => P_HR_NS239 <= P_HR_NS239 + T_N_STRESS;
                when "00101001100" => P_HR_NS240 <= P_HR_NS240 + T_N_STRESS;
                when "00101001110" => P_HR_NS241 <= P_HR_NS241 + T_N_STRESS;
                when "00101001111" => P_HR_NS242 <= P_HR_NS242 + T_N_STRESS;
                when "00101010000" => P_HR_NS243 <= P_HR_NS243 + T_N_STRESS;
                when "00101010001" => P_HR_NS244 <= P_HR_NS244 + T_N_STRESS;
                when "00101010010" => P_HR_NS245 <= P_HR_NS245 + T_N_STRESS;
                when "00101010011" => P_HR_NS246 <= P_HR_NS246 + T_N_STRESS;
                when "00101010100" => P_HR_NS247 <= P_HR_NS247 + T_N_STRESS;
                when "00101010101" => P_HR_NS248 <= P_HR_NS248 + T_N_STRESS;
                when "00101010110" => P_HR_NS249 <= P_HR_NS249 + T_N_STRESS;
                when "00101010111" => P_HR_NS250 <= P_HR_NS250 + T_N_STRESS;
                when "00101011000" => P_HR_NS251 <= P_HR_NS251 + T_N_STRESS;
                when "00101011001" => P_HR_NS252 <= P_HR_NS252 + T_N_STRESS;
                when "00101011010" => P_HR_NS253 <= P_HR_NS253 + T_N_STRESS;
                when "00101011011" => P_HR_NS254 <= P_HR_NS254 + T_N_STRESS;
                when "00101011100" => P_HR_NS255 <= P_HR_NS255 + T_N_STRESS;
                when "00101011101" => P_HR_NS256 <= P_HR_NS256 + T_N_STRESS;
                when "00101011110" => P_HR_NS257 <= P_HR_NS257 + T_N_STRESS;
                when "00101011111" => P_HR_NS258 <= P_HR_NS258 + T_N_STRESS;
                when "00101100000" => P_HR_NS259 <= P_HR_NS259 + T_N_STRESS;
                when "00101100001" => P_HR_NS260 <= P_HR_NS260 + T_N_STRESS;
                when "00101100010" => P_HR_NS261 <= P_HR_NS261 + T_N_STRESS;
                when "00101100011" => P_HR_NS262 <= P_HR_NS262 + T_N_STRESS;
                when "00101100100" => P_HR_NS263 <= P_HR_NS263 + T_N_STRESS;
                when "00101100101" => P_HR_NS264 <= P_HR_NS264 + T_N_STRESS;
                when "00101100110" => P_HR_NS265 <= P_HR_NS265 + T_N_STRESS;
                when "00101100111" => P_HR_NS266 <= P_HR_NS266 + T_N_STRESS;
                when "00101101000" => P_HR_NS267 <= P_HR_NS267 + T_N_STRESS;
                when "00101101001" => P_HR_NS268 <= P_HR_NS268 + T_N_STRESS;
                when "00101101010" => P_HR_NS269 <= P_HR_NS269 + T_N_STRESS;
                when "00101101011" => P_HR_NS270 <= P_HR_NS270 + T_N_STRESS;
                when "00101101100" => P_HR_NS271 <= P_HR_NS271 + T_N_STRESS;
                when "00101101101" => P_HR_NS272 <= P_HR_NS272 + T_N_STRESS;
                when "00101101110" => P_HR_NS273 <= P_HR_NS273 + T_N_STRESS;
                when "00101101111" => P_HR_NS274 <= P_HR_NS274 + T_N_STRESS;
                when "00101110000" => P_HR_NS275 <= P_HR_NS275 + T_N_STRESS;
                when "00101110001" => P_HR_NS276 <= P_HR_NS276 + T_N_STRESS;
                when "00101110010" => P_HR_NS277 <= P_HR_NS277 + T_N_STRESS;
                when "00101110011" => P_HR_NS278 <= P_HR_NS278 + T_N_STRESS;
                when "00101110100" => P_HR_NS279 <= P_HR_NS279 + T_N_STRESS;
                when "00101110101" => P_HR_NS280 <= P_HR_NS280 + T_N_STRESS;
                when "00101110110" => P_HR_NS281 <= P_HR_NS281 + T_N_STRESS;
                when "00101110111" => P_HR_NS282 <= P_HR_NS282 + T_N_STRESS;
                when "00101111000" => P_HR_NS283 <= P_HR_NS283 + T_N_STRESS;
                when "00101111001" => P_HR_NS284 <= P_HR_NS284 + T_N_STRESS;
                when "00101111010" => P_HR_NS285 <= P_HR_NS285 + T_N_STRESS;
                when "00101111011" => P_HR_NS286 <= P_HR_NS286 + T_N_STRESS;
                when "00101111100" => P_HR_NS287 <= P_HR_NS287 + T_N_STRESS;
                when "00101111101" => P_HR_NS288 <= P_HR_NS288 + T_N_STRESS;
                when "00101111110" => P_HR_NS289 <= P_HR_NS289 + T_N_STRESS;
                when "00101111111" => P_HR_NS290 <= P_HR_NS290 + T_N_STRESS;
                when "00110000000" => P_HR_NS291 <= P_HR_NS291 + T_N_STRESS;
                when "00110000001" => P_HR_NS292 <= P_HR_NS292 + T_N_STRESS;
                when "00110000010" => P_HR_NS293 <= P_HR_NS293 + T_N_STRESS;
                when "00110000011" => P_HR_NS294 <= P_HR_NS294 + T_N_STRESS;
                when "00110000100" => P_HR_NS295 <= P_HR_NS295 + T_N_STRESS;
                when "00110000101" => P_HR_NS296 <= P_HR_NS296 + T_N_STRESS;
                when "00110000110" => P_HR_NS297 <= P_HR_NS297 + T_N_STRESS;
                when "00110000111" => P_HR_NS298 <= P_HR_NS298 + T_N_STRESS;
                when "00110001000" => P_HR_NS299 <= P_HR_NS299 + T_N_STRESS;
                when "00110001001" => P_HR_NS300 <= P_HR_NS300 + T_N_STRESS;
                when "00110001010" => P_HR_NS301 <= P_HR_NS301 + T_N_STRESS;
                when "00110001011" => P_HR_NS302 <= P_HR_NS302 + T_N_STRESS;
                when "00110001100" => P_HR_NS303 <= P_HR_NS303 + T_N_STRESS;
                when "00110001101" => P_HR_NS304 <= P_HR_NS304 + T_N_STRESS;
                when "00110001110" => P_HR_NS305 <= P_HR_NS305 + T_N_STRESS;
                when "00110001111" => P_HR_NS306 <= P_HR_NS306 + T_N_STRESS;
                when "00110010000" => P_HR_NS307 <= P_HR_NS307 + T_N_STRESS;
                when "00110010001" => P_HR_NS308 <= P_HR_NS308 + T_N_STRESS;
                when "00110010010" => P_HR_NS309 <= P_HR_NS309 + T_N_STRESS;
                when "00110010011" => P_HR_NS310 <= P_HR_NS310 + T_N_STRESS;
                when "00110010100" => P_HR_NS311 <= P_HR_NS311 + T_N_STRESS;
                when "00110010101" => P_HR_NS312 <= P_HR_NS312 + T_N_STRESS;
                when "00110010110" => P_HR_NS313 <= P_HR_NS313 + T_N_STRESS;
                when "00110010111" => P_HR_NS314 <= P_HR_NS314 + T_N_STRESS;
                when "00110011000" => P_HR_NS315 <= P_HR_NS315 + T_N_STRESS;
                when "00110011001" => P_HR_NS316 <= P_HR_NS316 + T_N_STRESS;
                when "00110011010" => P_HR_NS317 <= P_HR_NS317 + T_N_STRESS;
                when "00110011011" => P_HR_NS318 <= P_HR_NS318 + T_N_STRESS;
                when "00110011100" => P_HR_NS319 <= P_HR_NS319 + T_N_STRESS;
                when "00110011101" => P_HR_NS320 <= P_HR_NS320 + T_N_STRESS;
                when "00110011110" => P_HR_NS321 <= P_HR_NS321 + T_N_STRESS;
                when "00110011111" => P_HR_NS322 <= P_HR_NS322 + T_N_STRESS;
                when "00110100000" => P_HR_NS323 <= P_HR_NS323 + T_N_STRESS;
                when "00110100001" => P_HR_NS324 <= P_HR_NS324 + T_N_STRESS;
                when "00110100010" => P_HR_NS325 <= P_HR_NS325 + T_N_STRESS;
                when "00110100011" => P_HR_NS326 <= P_HR_NS326 + T_N_STRESS;
                when "00110100100" => P_HR_NS327 <= P_HR_NS327 + T_N_STRESS;
                when "00110100101" => P_HR_NS328 <= P_HR_NS328 + T_N_STRESS;
                when "00110100110" => P_HR_NS329 <= P_HR_NS329 + T_N_STRESS;
                when "00110100111" => P_HR_NS330 <= P_HR_NS330 + T_N_STRESS;
                when "00110101000" => P_HR_NS331 <= P_HR_NS331 + T_N_STRESS;
                when "00110101001" => P_HR_NS332 <= P_HR_NS332 + T_N_STRESS;
                when "00110101010" => P_HR_NS333 <= P_HR_NS333 + T_N_STRESS;
                when "00110101011" => P_HR_NS334 <= P_HR_NS334 + T_N_STRESS;
                when "00110101100" => P_HR_NS335 <= P_HR_NS335 + T_N_STRESS;
                when "00110101101" => P_HR_NS336 <= P_HR_NS336 + T_N_STRESS;
                when "00110101110" => P_HR_NS337 <= P_HR_NS337 + T_N_STRESS;
                when "00110101111" => P_HR_NS338 <= P_HR_NS338 + T_N_STRESS;
                when "00110110000" => P_HR_NS339 <= P_HR_NS339 + T_N_STRESS;
                when "00110110001" => P_HR_NS340 <= P_HR_NS340 + T_N_STRESS;
                when "00110110010" => P_HR_NS341 <= P_HR_NS341 + T_N_STRESS;
                when "00110110011" => P_HR_NS342 <= P_HR_NS342 + T_N_STRESS;
                when "00110110100" => P_HR_NS343 <= P_HR_NS343 + T_N_STRESS;
                when "00110110101" => P_HR_NS344 <= P_HR_NS344 + T_N_STRESS;
                when "00110110110" => P_HR_NS345 <= P_HR_NS345 + T_N_STRESS;
                when "00110110111" => P_HR_NS346 <= P_HR_NS346 + T_N_STRESS;
                when "00110111000" => P_HR_NS347 <= P_HR_NS347 + T_N_STRESS;
                when "00110111001" => P_HR_NS348 <= P_HR_NS348 + T_N_STRESS;
                when "00110111010" => P_HR_NS349 <= P_HR_NS349 + T_N_STRESS;
                when "00110111011" => P_HR_NS350 <= P_HR_NS350 + T_N_STRESS;
                when "00110111100" => P_HR_NS351 <= P_HR_NS351 + T_N_STRESS;
                when "00110111101" => P_HR_NS352 <= P_HR_NS352 + T_N_STRESS;
                when "00110111110" => P_HR_NS353 <= P_HR_NS353 + T_N_STRESS;
                when "00110111111" => P_HR_NS354 <= P_HR_NS354 + T_N_STRESS;
                when "00111000000" => P_HR_NS355 <= P_HR_NS355 + T_N_STRESS;
                when "00111000001" => P_HR_NS356 <= P_HR_NS356 + T_N_STRESS;
                when "00111000010" => P_HR_NS357 <= P_HR_NS357 + T_N_STRESS;
                when "00111000011" => P_HR_NS358 <= P_HR_NS358 + T_N_STRESS;
                when "00111000100" => P_HR_NS359 <= P_HR_NS359 + T_N_STRESS;
                when "00111000101" => P_HR_NS360 <= P_HR_NS360 + T_N_STRESS;
                when "00111000110" => P_HR_NS361 <= P_HR_NS361 + T_N_STRESS;
                when "00111000111" => P_HR_NS362 <= P_HR_NS362 + T_N_STRESS;
                when "00111001000" => P_HR_NS363 <= P_HR_NS363 + T_N_STRESS;
                when "00111001001" => P_HR_NS364 <= P_HR_NS364 + T_N_STRESS;
                when "00111001010" => P_HR_NS365 <= P_HR_NS365 + T_N_STRESS;
                when "00111001011" => P_HR_NS366 <= P_HR_NS366 + T_N_STRESS;
                when "00111001100" => P_HR_NS367 <= P_HR_NS367 + T_N_STRESS;
                when "00111001101" => P_HR_NS368 <= P_HR_NS368 + T_N_STRESS;
                when "00111001110" => P_HR_NS369 <= P_HR_NS369 + T_N_STRESS;
                when "00111001111" => P_HR_NS370 <= P_HR_NS370 + T_N_STRESS;
                when "00111010000" => P_HR_NS371 <= P_HR_NS371 + T_N_STRESS;
                when "00111010001" => P_HR_NS372 <= P_HR_NS372 + T_N_STRESS;
                when "00111010010" => P_HR_NS373 <= P_HR_NS373 + T_N_STRESS;
                when "00111010011" => P_HR_NS374 <= P_HR_NS374 + T_N_STRESS;
                when "00111010100" => P_HR_NS375 <= P_HR_NS375 + T_N_STRESS;
                when "00111010101" => P_HR_NS376 <= P_HR_NS376 + T_N_STRESS;
                when "00111010110" => P_HR_NS377 <= P_HR_NS377 + T_N_STRESS;
                when "00111010111" => P_HR_NS378 <= P_HR_NS378 + T_N_STRESS;
                when "00111011000" => P_HR_NS379 <= P_HR_NS379 + T_N_STRESS;
                when "00111011001" => P_HR_NS380 <= P_HR_NS380 + T_N_STRESS;
                when "00111011010" => P_HR_NS381 <= P_HR_NS381 + T_N_STRESS;
                when "00111011011" => P_HR_NS382 <= P_HR_NS382 + T_N_STRESS;
                when "00111011100" => P_HR_NS383 <= P_HR_NS383 + T_N_STRESS;
                when "00111011101" => P_HR_NS384 <= P_HR_NS384 + T_N_STRESS;
                when "00111011110" => P_HR_NS385 <= P_HR_NS385 + T_N_STRESS;
                when "00111011111" => P_HR_NS386 <= P_HR_NS386 + T_N_STRESS;
                when "00111100000" => P_HR_NS387 <= P_HR_NS387 + T_N_STRESS;
                when "00111100001" => P_HR_NS388 <= P_HR_NS388 + T_N_STRESS;
                when "00111100010" => P_HR_NS389 <= P_HR_NS389 + T_N_STRESS;
                when "00111100011" => P_HR_NS390 <= P_HR_NS390 + T_N_STRESS;
                when "00111100100" => P_HR_NS391 <= P_HR_NS391 + T_N_STRESS;
                when "00111100101" => P_HR_NS392 <= P_HR_NS392 + T_N_STRESS;
                when "00111100110" => P_HR_NS393 <= P_HR_NS393 + T_N_STRESS;
                when "00111100111" => P_HR_NS394 <= P_HR_NS394 + T_N_STRESS;
                when "00111101000" => P_HR_NS395 <= P_HR_NS395 + T_N_STRESS;
                when "00111101001" => P_HR_NS396 <= P_HR_NS396 + T_N_STRESS;
                when "00111101010" => P_HR_NS397 <= P_HR_NS397 + T_N_STRESS;
                when "00111101011" => P_HR_NS398 <= P_HR_NS398 + T_N_STRESS;
                when "00111101100" => P_HR_NS399 <= P_HR_NS399 + T_N_STRESS;
                when "00111101101" => P_HR_NS400 <= P_HR_NS400 + T_N_STRESS;
                when "00111101110" => P_HR_NS401 <= P_HR_NS401 + T_N_STRESS;
                when "00111101111" => P_HR_NS402 <= P_HR_NS402 + T_N_STRESS;
                when "00111110000" => P_HR_NS403 <= P_HR_NS403 + T_N_STRESS;
                when "00111110001" => P_HR_NS404 <= P_HR_NS404 + T_N_STRESS;
                when "00111110010" => P_HR_NS405 <= P_HR_NS405 + T_N_STRESS;
                when "00111110011" => P_HR_NS406 <= P_HR_NS406 + T_N_STRESS;
                when "00111110100" => P_HR_NS407 <= P_HR_NS407 + T_N_STRESS;
                when "00111110101" => P_HR_NS408 <= P_HR_NS408 + T_N_STRESS;
                when "00111110110" => P_HR_NS409 <= P_HR_NS409 + T_N_STRESS;
                when "00111110111" => P_HR_NS410 <= P_HR_NS410 + T_N_STRESS;
                when "00111111000" => P_HR_NS411 <= P_HR_NS411 + T_N_STRESS;
                when "00111111001" => P_HR_NS412 <= P_HR_NS412 + T_N_STRESS;
                when "00111111010" => P_HR_NS413 <= P_HR_NS413 + T_N_STRESS;
                when "00111111011" => P_HR_NS414 <= P_HR_NS414 + T_N_STRESS;
                when "00111111100" => P_HR_NS415 <= P_HR_NS415 + T_N_STRESS;
                when "00111111101" => P_HR_NS416 <= P_HR_NS416 + T_N_STRESS;
                when "00111111110" => P_HR_NS417 <= P_HR_NS417 + T_N_STRESS;
                when "00111111111" => P_HR_NS418 <= P_HR_NS418 + T_N_STRESS;
                when "01000000000" => P_HR_NS419 <= P_HR_NS419 + T_N_STRESS;
                when "01000000001" => P_HR_NS420 <= P_HR_NS420 + T_N_STRESS;
                when "01000000010" => P_HR_NS421 <= P_HR_NS421 + T_N_STRESS;
                when "01000000011" => P_HR_NS422 <= P_HR_NS422 + T_N_STRESS;
                when "01000000100" => P_HR_NS423 <= P_HR_NS423 + T_N_STRESS;
                when "01000000101" => P_HR_NS424 <= P_HR_NS424 + T_N_STRESS;
                when "01000000110" => P_HR_NS425 <= P_HR_NS425 + T_N_STRESS;
                when "01000000111" => P_HR_NS426 <= P_HR_NS426 + T_N_STRESS;
                when "01000001000" => P_HR_NS427 <= P_HR_NS427 + T_N_STRESS;
                when "01000001001" => P_HR_NS428 <= P_HR_NS428 + T_N_STRESS;
                when "01000001010" => P_HR_NS429 <= P_HR_NS429 + T_N_STRESS;
                when "01000001011" => P_HR_NS430 <= P_HR_NS430 + T_N_STRESS;
                when "01000001100" => P_HR_NS431 <= P_HR_NS431 + T_N_STRESS;
                when "01000001101" => P_HR_NS432 <= P_HR_NS432 + T_N_STRESS;
                when "01000001110" => P_HR_NS433 <= P_HR_NS433 + T_N_STRESS;
                when "01000001111" => P_HR_NS434 <= P_HR_NS434 + T_N_STRESS;
                when "01000010000" => P_HR_NS435 <= P_HR_NS435 + T_N_STRESS;
                when "01000010001" => P_HR_NS436 <= P_HR_NS436 + T_N_STRESS;
                when "01000010010" => P_HR_NS437 <= P_HR_NS437 + T_N_STRESS;
                when "01000010011" => P_HR_NS438 <= P_HR_NS438 + T_N_STRESS;
                when "01000010100" => P_HR_NS439 <= P_HR_NS439 + T_N_STRESS;
                when "01000010101" => P_HR_NS440 <= P_HR_NS440 + T_N_STRESS;
                when "01000010110" => P_HR_NS441 <= P_HR_NS441 + T_N_STRESS;
                when "01000010111" => P_HR_NS442 <= P_HR_NS442 + T_N_STRESS;
                when "01000011000" => P_HR_NS443 <= P_HR_NS443 + T_N_STRESS;
                when "01000011001" => P_HR_NS444 <= P_HR_NS444 + T_N_STRESS;
                when "01000011010" => P_HR_NS445 <= P_HR_NS445 + T_N_STRESS;
                when "01000011011" => P_HR_NS446 <= P_HR_NS446 + T_N_STRESS;
                when "01000011100" => P_HR_NS447 <= P_HR_NS447 + T_N_STRESS;
                when "01000011101" => P_HR_NS448 <= P_HR_NS448 + T_N_STRESS;
                when "01000011110" => P_HR_NS449 <= P_HR_NS449 + T_N_STRESS;
                when "01000011111" => P_HR_NS450 <= P_HR_NS450 + T_N_STRESS;
                when "01000100000" => P_HR_NS451 <= P_HR_NS451 + T_N_STRESS;
                when "01000100001" => P_HR_NS452 <= P_HR_NS452 + T_N_STRESS;
                when "01000100010" => P_HR_NS453 <= P_HR_NS453 + T_N_STRESS;
                when "01000100011" => P_HR_NS454 <= P_HR_NS454 + T_N_STRESS;
                when "01000100100" => P_HR_NS455 <= P_HR_NS455 + T_N_STRESS;
                when "01000100101" => P_HR_NS456 <= P_HR_NS456 + T_N_STRESS;
                when "01000100110" => P_HR_NS457 <= P_HR_NS457 + T_N_STRESS;
                when "01000100111" => P_HR_NS458 <= P_HR_NS458 + T_N_STRESS;
                when "01000101000" => P_HR_NS459 <= P_HR_NS459 + T_N_STRESS;
                when "01000101001" => P_HR_NS460 <= P_HR_NS460 + T_N_STRESS;
                when "01000101010" => P_HR_NS461 <= P_HR_NS461 + T_N_STRESS;
                when "01000101011" => P_HR_NS462 <= P_HR_NS462 + T_N_STRESS;
                when "01000101100" => P_HR_NS463 <= P_HR_NS463 + T_N_STRESS;
                when "01000101101" => P_HR_NS464 <= P_HR_NS464 + T_N_STRESS;
                when "01000101110" => P_HR_NS465 <= P_HR_NS465 + T_N_STRESS;
                when "01000101111" => P_HR_NS466 <= P_HR_NS466 + T_N_STRESS;
                when "01000110000" => P_HR_NS467 <= P_HR_NS467 + T_N_STRESS;
                when "01000110001" => P_HR_NS468 <= P_HR_NS468 + T_N_STRESS;
                when "01000110010" => P_HR_NS469 <= P_HR_NS469 + T_N_STRESS;
                when "01000110011" => P_HR_NS470 <= P_HR_NS470 + T_N_STRESS;
                when "01000110100" => P_HR_NS471 <= P_HR_NS471 + T_N_STRESS;
                when "01000110101" => P_HR_NS472 <= P_HR_NS472 + T_N_STRESS;
                when "01000110110" => P_HR_NS473 <= P_HR_NS473 + T_N_STRESS;
                when "01000110111" => P_HR_NS474 <= P_HR_NS474 + T_N_STRESS;
                when "01000111000" => P_HR_NS475 <= P_HR_NS475 + T_N_STRESS;
                when "01000111001" => P_HR_NS476 <= P_HR_NS476 + T_N_STRESS;
                when "01000111010" => P_HR_NS477 <= P_HR_NS477 + T_N_STRESS;
                when "01000111011" => P_HR_NS478 <= P_HR_NS478 + T_N_STRESS;
                when "01000111100" => P_HR_NS479 <= P_HR_NS479 + T_N_STRESS;
                when "01000111101" => P_HR_NS480 <= P_HR_NS480 + T_N_STRESS;
                when "01000111110" => P_HR_NS481 <= P_HR_NS481 + T_N_STRESS;
                when "01000111111" => P_HR_NS482 <= P_HR_NS482 + T_N_STRESS;
                when "01001000000" => P_HR_NS483 <= P_HR_NS483 + T_N_STRESS;
                when "01001000001" => P_HR_NS484 <= P_HR_NS484 + T_N_STRESS;
                when "01001000010" => P_HR_NS485 <= P_HR_NS485 + T_N_STRESS;
                when "01001000011" => P_HR_NS486 <= P_HR_NS486 + T_N_STRESS;
                when "01001000100" => P_HR_NS487 <= P_HR_NS487 + T_N_STRESS;
                when "01001000101" => P_HR_NS488 <= P_HR_NS488 + T_N_STRESS;
                when "01001000110" => P_HR_NS489 <= P_HR_NS489 + T_N_STRESS;
                when "01001000111" => P_HR_NS490 <= P_HR_NS490 + T_N_STRESS;
                when "01001001000" => P_HR_NS491 <= P_HR_NS491 + T_N_STRESS;
                when "01001001001" => P_HR_NS492 <= P_HR_NS492 + T_N_STRESS;
                when "01001001010" => P_HR_NS493 <= P_HR_NS493 + T_N_STRESS;
                when "01001001011" => P_HR_NS494 <= P_HR_NS494 + T_N_STRESS;
                when "01001001100" => P_HR_NS495 <= P_HR_NS495 + T_N_STRESS;
                when "01001001101" => P_HR_NS496 <= P_HR_NS496 + T_N_STRESS;
                when "01001001111" => P_HR_NS497 <= P_HR_NS497 + T_N_STRESS;
                when "01001010000" => P_HR_NS498 <= P_HR_NS498 + T_N_STRESS;
                when "01001010001" => P_HR_NS499 <= P_HR_NS499 + T_N_STRESS;
                when "01001010010" => P_HR_NS500 <= P_HR_NS500 + T_N_STRESS;
                when "01001010011" => P_HR_NS501 <= P_HR_NS501 + T_N_STRESS;
                when "01001010100" => P_HR_NS502 <= P_HR_NS502 + T_N_STRESS;
                when "01001010101" => P_HR_NS503 <= P_HR_NS503 + T_N_STRESS;
                when "01001010110" => P_HR_NS504 <= P_HR_NS504 + T_N_STRESS;
                when "01001010111" => P_HR_NS505 <= P_HR_NS505 + T_N_STRESS;
                when "01001011000" => P_HR_NS506 <= P_HR_NS506 + T_N_STRESS;
                when "01001011001" => P_HR_NS507 <= P_HR_NS507 + T_N_STRESS;
                when "01001011010" => P_HR_NS508 <= P_HR_NS508 + T_N_STRESS;
                when "01001011011" => P_HR_NS509 <= P_HR_NS509 + T_N_STRESS;
                when "01001011100" => P_HR_NS510 <= P_HR_NS510 + T_N_STRESS;
                when "01001011101" => P_HR_NS511 <= P_HR_NS511 + T_N_STRESS;
                when "01001011110" => P_HR_NS512 <= P_HR_NS512 + T_N_STRESS;
                when "01001100000" => P_HR_NS513 <= P_HR_NS513 + T_N_STRESS;
                when "01001100001" => P_HR_NS514 <= P_HR_NS514 + T_N_STRESS;
                when "01001100010" => P_HR_NS515 <= P_HR_NS515 + T_N_STRESS;
                when "01001100011" => P_HR_NS516 <= P_HR_NS516 + T_N_STRESS;
                when "01001100100" => P_HR_NS517 <= P_HR_NS517 + T_N_STRESS;
                when "01001100101" => P_HR_NS518 <= P_HR_NS518 + T_N_STRESS;
                when "01001100110" => P_HR_NS519 <= P_HR_NS519 + T_N_STRESS;
                when "01001100111" => P_HR_NS520 <= P_HR_NS520 + T_N_STRESS;
                when "01001101001" => P_HR_NS521 <= P_HR_NS521 + T_N_STRESS;
                when "01001101010" => P_HR_NS522 <= P_HR_NS522 + T_N_STRESS;
                when "01001101011" => P_HR_NS523 <= P_HR_NS523 + T_N_STRESS;
                when "01001101100" => P_HR_NS524 <= P_HR_NS524 + T_N_STRESS;
                when "01001101101" => P_HR_NS525 <= P_HR_NS525 + T_N_STRESS;
                when "01001101110" => P_HR_NS526 <= P_HR_NS526 + T_N_STRESS;
                when "01001101111" => P_HR_NS527 <= P_HR_NS527 + T_N_STRESS;
                when "01001110001" => P_HR_NS528 <= P_HR_NS528 + T_N_STRESS;
                when "01001110010" => P_HR_NS529 <= P_HR_NS529 + T_N_STRESS;
                when "01001110011" => P_HR_NS530 <= P_HR_NS530 + T_N_STRESS;
                when "01001110100" => P_HR_NS531 <= P_HR_NS531 + T_N_STRESS;
                when "01001110101" => P_HR_NS532 <= P_HR_NS532 + T_N_STRESS;
                when "01001110110" => P_HR_NS533 <= P_HR_NS533 + T_N_STRESS;
                when "01001111000" => P_HR_NS534 <= P_HR_NS534 + T_N_STRESS;
                when "01001111001" => P_HR_NS535 <= P_HR_NS535 + T_N_STRESS;
                when "01001111010" => P_HR_NS536 <= P_HR_NS536 + T_N_STRESS;
                when "01001111011" => P_HR_NS537 <= P_HR_NS537 + T_N_STRESS;
                when "01001111100" => P_HR_NS538 <= P_HR_NS538 + T_N_STRESS;
                when "01001111110" => P_HR_NS539 <= P_HR_NS539 + T_N_STRESS;
                when "01001111111" => P_HR_NS540 <= P_HR_NS540 + T_N_STRESS;
                when "01010000000" => P_HR_NS541 <= P_HR_NS541 + T_N_STRESS;
                when "01010000001" => P_HR_NS542 <= P_HR_NS542 + T_N_STRESS;
                when "01010000010" => P_HR_NS543 <= P_HR_NS543 + T_N_STRESS;
                when "01010000100" => P_HR_NS544 <= P_HR_NS544 + T_N_STRESS;
                when "01010000101" => P_HR_NS545 <= P_HR_NS545 + T_N_STRESS;
                when "01010000110" => P_HR_NS546 <= P_HR_NS546 + T_N_STRESS;
                when "01010000111" => P_HR_NS547 <= P_HR_NS547 + T_N_STRESS;
                when "01010001001" => P_HR_NS548 <= P_HR_NS548 + T_N_STRESS;
                when "01010001010" => P_HR_NS549 <= P_HR_NS549 + T_N_STRESS;
                when "01010001011" => P_HR_NS550 <= P_HR_NS550 + T_N_STRESS;
                when "01010001100" => P_HR_NS551 <= P_HR_NS551 + T_N_STRESS;
                when "01010001110" => P_HR_NS552 <= P_HR_NS552 + T_N_STRESS;
                when "01010001111" => P_HR_NS553 <= P_HR_NS553 + T_N_STRESS;
                when "01010010000" => P_HR_NS554 <= P_HR_NS554 + T_N_STRESS;
                when "01010010010" => P_HR_NS555 <= P_HR_NS555 + T_N_STRESS;
                when "01010010011" => P_HR_NS556 <= P_HR_NS556 + T_N_STRESS;
                when "01010010100" => P_HR_NS557 <= P_HR_NS557 + T_N_STRESS;
                when "01010010101" => P_HR_NS558 <= P_HR_NS558 + T_N_STRESS;
                when "01010010111" => P_HR_NS559 <= P_HR_NS559 + T_N_STRESS;
                when "01010011000" => P_HR_NS560 <= P_HR_NS560 + T_N_STRESS;
                when "01010011001" => P_HR_NS561 <= P_HR_NS561 + T_N_STRESS;
                when "01010011011" => P_HR_NS562 <= P_HR_NS562 + T_N_STRESS;
                when "01010011100" => P_HR_NS563 <= P_HR_NS563 + T_N_STRESS;
                when "01010011101" => P_HR_NS564 <= P_HR_NS564 + T_N_STRESS;
                when "01010011111" => P_HR_NS565 <= P_HR_NS565 + T_N_STRESS;
                when "01010100000" => P_HR_NS566 <= P_HR_NS566 + T_N_STRESS;
                when "01010100001" => P_HR_NS567 <= P_HR_NS567 + T_N_STRESS;
                when "01010100011" => P_HR_NS568 <= P_HR_NS568 + T_N_STRESS;
                when "01010100100" => P_HR_NS569 <= P_HR_NS569 + T_N_STRESS;
                when "01010100101" => P_HR_NS570 <= P_HR_NS570 + T_N_STRESS;
                when "01010100111" => P_HR_NS571 <= P_HR_NS571 + T_N_STRESS;
                when "01010101000" => P_HR_NS572 <= P_HR_NS572 + T_N_STRESS;
                when "01010101010" => P_HR_NS573 <= P_HR_NS573 + T_N_STRESS;
                when "01010101011" => P_HR_NS574 <= P_HR_NS574 + T_N_STRESS;
                when "01010101100" => P_HR_NS575 <= P_HR_NS575 + T_N_STRESS;
                when "01010101110" => P_HR_NS576 <= P_HR_NS576 + T_N_STRESS;
                when "01010101111" => P_HR_NS577 <= P_HR_NS577 + T_N_STRESS;
                when "01010110001" => P_HR_NS578 <= P_HR_NS578 + T_N_STRESS;
                when "01010110010" => P_HR_NS579 <= P_HR_NS579 + T_N_STRESS;
                when "01010110011" => P_HR_NS580 <= P_HR_NS580 + T_N_STRESS;
                when "01010110101" => P_HR_NS581 <= P_HR_NS581 + T_N_STRESS;
                when "01010110110" => P_HR_NS582 <= P_HR_NS582 + T_N_STRESS;
                when "01010111000" => P_HR_NS583 <= P_HR_NS583 + T_N_STRESS;
                when "01010111001" => P_HR_NS584 <= P_HR_NS584 + T_N_STRESS;
                when "01010111011" => P_HR_NS585 <= P_HR_NS585 + T_N_STRESS;
                when "01010111100" => P_HR_NS586 <= P_HR_NS586 + T_N_STRESS;
                when "01010111101" => P_HR_NS587 <= P_HR_NS587 + T_N_STRESS;
                when "01010111111" => P_HR_NS588 <= P_HR_NS588 + T_N_STRESS;
                when "01011000000" => P_HR_NS589 <= P_HR_NS589 + T_N_STRESS;
                when "01011000010" => P_HR_NS590 <= P_HR_NS590 + T_N_STRESS;
                when "01011000011" => P_HR_NS591 <= P_HR_NS591 + T_N_STRESS;
                when "01011000101" => P_HR_NS592 <= P_HR_NS592 + T_N_STRESS;
                when "01011000110" => P_HR_NS593 <= P_HR_NS593 + T_N_STRESS;
                when "01011001000" => P_HR_NS594 <= P_HR_NS594 + T_N_STRESS;
                when "01011001001" => P_HR_NS595 <= P_HR_NS595 + T_N_STRESS;
                when "01011001011" => P_HR_NS596 <= P_HR_NS596 + T_N_STRESS;
                when "01011001100" => P_HR_NS597 <= P_HR_NS597 + T_N_STRESS;
                when "01011001110" => P_HR_NS598 <= P_HR_NS598 + T_N_STRESS;
                when "01011001111" => P_HR_NS599 <= P_HR_NS599 + T_N_STRESS;
                when "01011010001" => P_HR_NS600 <= P_HR_NS600 + T_N_STRESS;
                when "01011010011" => P_HR_NS601 <= P_HR_NS601 + T_N_STRESS;
                when "01011010100" => P_HR_NS602 <= P_HR_NS602 + T_N_STRESS;
                when "01011010110" => P_HR_NS603 <= P_HR_NS603 + T_N_STRESS;
                when "01011010111" => P_HR_NS604 <= P_HR_NS604 + T_N_STRESS;
                when "01011011001" => P_HR_NS605 <= P_HR_NS605 + T_N_STRESS;
                when "01011011010" => P_HR_NS606 <= P_HR_NS606 + T_N_STRESS;
                when "01011011100" => P_HR_NS607 <= P_HR_NS607 + T_N_STRESS;
                when "01011011110" => P_HR_NS608 <= P_HR_NS608 + T_N_STRESS;
                when "01011011111" => P_HR_NS609 <= P_HR_NS609 + T_N_STRESS;
                when "01011100001" => P_HR_NS610 <= P_HR_NS610 + T_N_STRESS;
                when "01011100010" => P_HR_NS611 <= P_HR_NS611 + T_N_STRESS;
                when "01011100100" => P_HR_NS612 <= P_HR_NS612 + T_N_STRESS;
                when "01011100110" => P_HR_NS613 <= P_HR_NS613 + T_N_STRESS;
                when "01011100111" => P_HR_NS614 <= P_HR_NS614 + T_N_STRESS;
                when "01011101001" => P_HR_NS615 <= P_HR_NS615 + T_N_STRESS;
                when "01011101011" => P_HR_NS616 <= P_HR_NS616 + T_N_STRESS;
                when "01011101100" => P_HR_NS617 <= P_HR_NS617 + T_N_STRESS;
                when "01011101110" => P_HR_NS618 <= P_HR_NS618 + T_N_STRESS;
                when "01011110000" => P_HR_NS619 <= P_HR_NS619 + T_N_STRESS;
                when "01011110001" => P_HR_NS620 <= P_HR_NS620 + T_N_STRESS;
                when "01011110011" => P_HR_NS621 <= P_HR_NS621 + T_N_STRESS;
                when "01011110101" => P_HR_NS622 <= P_HR_NS622 + T_N_STRESS;
                when "01011110110" => P_HR_NS623 <= P_HR_NS623 + T_N_STRESS;
                when "01011111000" => P_HR_NS624 <= P_HR_NS624 + T_N_STRESS;
                when "01011111010" => P_HR_NS625 <= P_HR_NS625 + T_N_STRESS;
                when "01011111100" => P_HR_NS626 <= P_HR_NS626 + T_N_STRESS;
                when "01011111101" => P_HR_NS627 <= P_HR_NS627 + T_N_STRESS;
                when "01011111111" => P_HR_NS628 <= P_HR_NS628 + T_N_STRESS;
                when "01100000001" => P_HR_NS629 <= P_HR_NS629 + T_N_STRESS;
                when "01100000011" => P_HR_NS630 <= P_HR_NS630 + T_N_STRESS;
                when "01100000100" => P_HR_NS631 <= P_HR_NS631 + T_N_STRESS;
                when "01100000110" => P_HR_NS632 <= P_HR_NS632 + T_N_STRESS;
                when "01100001000" => P_HR_NS633 <= P_HR_NS633 + T_N_STRESS;
                when "01100001010" => P_HR_NS634 <= P_HR_NS634 + T_N_STRESS;
                when "01100001100" => P_HR_NS635 <= P_HR_NS635 + T_N_STRESS;
                when "01100001101" => P_HR_NS636 <= P_HR_NS636 + T_N_STRESS;
                when "01100001111" => P_HR_NS637 <= P_HR_NS637 + T_N_STRESS;
                when "01100010001" => P_HR_NS638 <= P_HR_NS638 + T_N_STRESS;
                when "01100010011" => P_HR_NS639 <= P_HR_NS639 + T_N_STRESS;
                when "01100010101" => P_HR_NS640 <= P_HR_NS640 + T_N_STRESS;
                when "01100010111" => P_HR_NS641 <= P_HR_NS641 + T_N_STRESS;
                when "01100011000" => P_HR_NS642 <= P_HR_NS642 + T_N_STRESS;
                when "01100011010" => P_HR_NS643 <= P_HR_NS643 + T_N_STRESS;
                when "01100011100" => P_HR_NS644 <= P_HR_NS644 + T_N_STRESS;
                when "01100011110" => P_HR_NS645 <= P_HR_NS645 + T_N_STRESS;
                when "01100100000" => P_HR_NS646 <= P_HR_NS646 + T_N_STRESS;
                when "01100100010" => P_HR_NS647 <= P_HR_NS647 + T_N_STRESS;
                when "01100100100" => P_HR_NS648 <= P_HR_NS648 + T_N_STRESS;
                when "01100100110" => P_HR_NS649 <= P_HR_NS649 + T_N_STRESS;
                when "01100101000" => P_HR_NS650 <= P_HR_NS650 + T_N_STRESS;
                when "01100101010" => P_HR_NS651 <= P_HR_NS651 + T_N_STRESS;
                when "01100101100" => P_HR_NS652 <= P_HR_NS652 + T_N_STRESS;
                when "01100101110" => P_HR_NS653 <= P_HR_NS653 + T_N_STRESS;
                when "01100110000" => P_HR_NS654 <= P_HR_NS654 + T_N_STRESS;
                when "01100110010" => P_HR_NS655 <= P_HR_NS655 + T_N_STRESS;
                when "01100110100" => P_HR_NS656 <= P_HR_NS656 + T_N_STRESS;
                when "01100110110" => P_HR_NS657 <= P_HR_NS657 + T_N_STRESS;
                when "01100111000" => P_HR_NS658 <= P_HR_NS658 + T_N_STRESS;
                when "01100111010" => P_HR_NS659 <= P_HR_NS659 + T_N_STRESS;
                when "01100111100" => P_HR_NS660 <= P_HR_NS660 + T_N_STRESS;
                when "01100111110" => P_HR_NS661 <= P_HR_NS661 + T_N_STRESS;
                when "01101000000" => P_HR_NS662 <= P_HR_NS662 + T_N_STRESS;
                when "01101000010" => P_HR_NS663 <= P_HR_NS663 + T_N_STRESS;
                when "01101000100" => P_HR_NS664 <= P_HR_NS664 + T_N_STRESS;
                when "01101000110" => P_HR_NS665 <= P_HR_NS665 + T_N_STRESS;
                when "01101001000" => P_HR_NS666 <= P_HR_NS666 + T_N_STRESS;
                when "01101001010" => P_HR_NS667 <= P_HR_NS667 + T_N_STRESS;
                when "01101001100" => P_HR_NS668 <= P_HR_NS668 + T_N_STRESS;
                when "01101001110" => P_HR_NS669 <= P_HR_NS669 + T_N_STRESS;
                when "01101010000" => P_HR_NS670 <= P_HR_NS670 + T_N_STRESS;
                when "01101010011" => P_HR_NS671 <= P_HR_NS671 + T_N_STRESS;
                when "01101010101" => P_HR_NS672 <= P_HR_NS672 + T_N_STRESS;
                when "01101010111" => P_HR_NS673 <= P_HR_NS673 + T_N_STRESS;
                when "01101011001" => P_HR_NS674 <= P_HR_NS674 + T_N_STRESS;
                when "01101011011" => P_HR_NS675 <= P_HR_NS675 + T_N_STRESS;
                when "01101011110" => P_HR_NS676 <= P_HR_NS676 + T_N_STRESS;
                when "01101100000" => P_HR_NS677 <= P_HR_NS677 + T_N_STRESS;
                when "01101100010" => P_HR_NS678 <= P_HR_NS678 + T_N_STRESS;
                when "01101100100" => P_HR_NS679 <= P_HR_NS679 + T_N_STRESS;
                when "01101100110" => P_HR_NS680 <= P_HR_NS680 + T_N_STRESS;
                when "01101101001" => P_HR_NS681 <= P_HR_NS681 + T_N_STRESS;
                when "01101101011" => P_HR_NS682 <= P_HR_NS682 + T_N_STRESS;
                when "01101101101" => P_HR_NS683 <= P_HR_NS683 + T_N_STRESS;
                when "01101110000" => P_HR_NS684 <= P_HR_NS684 + T_N_STRESS;
                when "01101110010" => P_HR_NS685 <= P_HR_NS685 + T_N_STRESS;
                when "01101110100" => P_HR_NS686 <= P_HR_NS686 + T_N_STRESS;
                when "01101110111" => P_HR_NS687 <= P_HR_NS687 + T_N_STRESS;
                when "01101111001" => P_HR_NS688 <= P_HR_NS688 + T_N_STRESS;
                when "01101111011" => P_HR_NS689 <= P_HR_NS689 + T_N_STRESS;
                when "01101111110" => P_HR_NS690 <= P_HR_NS690 + T_N_STRESS;
                when "01110000000" => P_HR_NS691 <= P_HR_NS691 + T_N_STRESS;
                when "01110000010" => P_HR_NS692 <= P_HR_NS692 + T_N_STRESS;
                when "01110000101" => P_HR_NS693 <= P_HR_NS693 + T_N_STRESS;
                when "01110000111" => P_HR_NS694 <= P_HR_NS694 + T_N_STRESS;
                when "01110001010" => P_HR_NS695 <= P_HR_NS695 + T_N_STRESS;
                when "01110001100" => P_HR_NS696 <= P_HR_NS696 + T_N_STRESS;
                when "01110001111" => P_HR_NS697 <= P_HR_NS697 + T_N_STRESS;
                when "01110010001" => P_HR_NS698 <= P_HR_NS698 + T_N_STRESS;
                when "01110010100" => P_HR_NS699 <= P_HR_NS699 + T_N_STRESS;
                when "01110010110" => P_HR_NS700 <= P_HR_NS700 + T_N_STRESS;
                when "01110011001" => P_HR_NS701 <= P_HR_NS701 + T_N_STRESS;
                when "01110011011" => P_HR_NS702 <= P_HR_NS702 + T_N_STRESS;
                when "01110011110" => P_HR_NS703 <= P_HR_NS703 + T_N_STRESS;
                when "01110100000" => P_HR_NS704 <= P_HR_NS704 + T_N_STRESS;
                when "01110100011" => P_HR_NS705 <= P_HR_NS705 + T_N_STRESS;
                when "01110101000" => P_HR_NS706 <= P_HR_NS706 + T_N_STRESS;
                when "01110101011" => P_HR_NS707 <= P_HR_NS707 + T_N_STRESS;
                when "01110101101" => P_HR_NS708 <= P_HR_NS708 + T_N_STRESS;
                when "01110110000" => P_HR_NS709 <= P_HR_NS709 + T_N_STRESS;
                when "01110110101" => P_HR_NS710 <= P_HR_NS710 + T_N_STRESS;
                when "01110111000" => P_HR_NS711 <= P_HR_NS711 + T_N_STRESS;
                when "01110111011" => P_HR_NS712 <= P_HR_NS712 + T_N_STRESS;
                when "01110111101" => P_HR_NS713 <= P_HR_NS713 + T_N_STRESS;
                when "01111001011" => P_HR_NS714 <= P_HR_NS714 + T_N_STRESS;
                when "01111010001" => P_HR_NS715 <= P_HR_NS715 + T_N_STRESS;
                when "01111011001" => P_HR_NS716 <= P_HR_NS716 + T_N_STRESS;
                when "01111011100" => P_HR_NS717 <= P_HR_NS717 + T_N_STRESS;
                when "01111100101" => P_HR_NS718 <= P_HR_NS718 + T_N_STRESS;
                when "10010000011" => P_HR_NS719 <= P_HR_NS719 + T_N_STRESS;
                when "10010011011" => P_HR_NS720 <= P_HR_NS720 + T_N_STRESS;
                when "10100101011" => P_HR_NS721 <= P_HR_NS721 + T_N_STRESS;
                when "10101100001" => P_HR_NS722 <= P_HR_NS722 + T_N_STRESS;
                when "10101100111" => P_HR_NS723 <= P_HR_NS723 + T_N_STRESS;
                when "10110011100" => P_HR_NS724 <= P_HR_NS724 + T_N_STRESS;
                when "11100000101" => P_HR_NS725 <= P_HR_NS725 + T_N_STRESS;
                when "11110101101" => P_HR_NS726 <= P_HR_NS726 + T_N_STRESS;
				when others            => null;
			end case;

			case eda is
                when "00000010" => P_EDA_NS1 <= P_EDA_NS1 + T_N_STRESS;
                when "00000011" => P_EDA_NS2 <= P_EDA_NS2 + T_N_STRESS;
                when "00000100" => P_EDA_NS3 <= P_EDA_NS3 + T_N_STRESS;
                when "00000101" => P_EDA_NS4 <= P_EDA_NS4 + T_N_STRESS;
                when "00000110" => P_EDA_NS5 <= P_EDA_NS5 + T_N_STRESS;
                when "00000111" => P_EDA_NS6 <= P_EDA_NS6 + T_N_STRESS;
                when "00001000" => P_EDA_NS7 <= P_EDA_NS7 + T_N_STRESS;
                when "00001001" => P_EDA_NS8 <= P_EDA_NS8 + T_N_STRESS;
                when "00001010" => P_EDA_NS9 <= P_EDA_NS9 + T_N_STRESS;
                when "00001011" => P_EDA_NS10 <= P_EDA_NS10 + T_N_STRESS;
                when "00001100" => P_EDA_NS11 <= P_EDA_NS11 + T_N_STRESS;
                when "00001101" => P_EDA_NS12 <= P_EDA_NS12 + T_N_STRESS;
                when "00001110" => P_EDA_NS13 <= P_EDA_NS13 + T_N_STRESS;
                when "00001111" => P_EDA_NS14 <= P_EDA_NS14 + T_N_STRESS;
                when "00010000" => P_EDA_NS15 <= P_EDA_NS15 + T_N_STRESS;
                when "00010001" => P_EDA_NS16 <= P_EDA_NS16 + T_N_STRESS;
                when "00010010" => P_EDA_NS17 <= P_EDA_NS17 + T_N_STRESS;
                when "00010011" => P_EDA_NS18 <= P_EDA_NS18 + T_N_STRESS;
                when "00010100" => P_EDA_NS19 <= P_EDA_NS19 + T_N_STRESS;
                when "00010101" => P_EDA_NS20 <= P_EDA_NS20 + T_N_STRESS;
                when "00010110" => P_EDA_NS21 <= P_EDA_NS21 + T_N_STRESS;
                when "00010111" => P_EDA_NS22 <= P_EDA_NS22 + T_N_STRESS;
                when "00011000" => P_EDA_NS23 <= P_EDA_NS23 + T_N_STRESS;
                when "00011001" => P_EDA_NS24 <= P_EDA_NS24 + T_N_STRESS;
                when "00011010" => P_EDA_NS25 <= P_EDA_NS25 + T_N_STRESS;
                when "00011011" => P_EDA_NS26 <= P_EDA_NS26 + T_N_STRESS;
                when "00011100" => P_EDA_NS27 <= P_EDA_NS27 + T_N_STRESS;
                when "00011101" => P_EDA_NS28 <= P_EDA_NS28 + T_N_STRESS;
                when "00011110" => P_EDA_NS29 <= P_EDA_NS29 + T_N_STRESS;
                when "00011111" => P_EDA_NS30 <= P_EDA_NS30 + T_N_STRESS;
                when "00100000" => P_EDA_NS31 <= P_EDA_NS31 + T_N_STRESS;
                when "00100001" => P_EDA_NS32 <= P_EDA_NS32 + T_N_STRESS;
                when "00100010" => P_EDA_NS33 <= P_EDA_NS33 + T_N_STRESS;
                when "00100011" => P_EDA_NS34 <= P_EDA_NS34 + T_N_STRESS;
                when "00100100" => P_EDA_NS35 <= P_EDA_NS35 + T_N_STRESS;
                when "00100101" => P_EDA_NS36 <= P_EDA_NS36 + T_N_STRESS;
                when "00100110" => P_EDA_NS37 <= P_EDA_NS37 + T_N_STRESS;
                when "00100111" => P_EDA_NS38 <= P_EDA_NS38 + T_N_STRESS;
                when "00101000" => P_EDA_NS39 <= P_EDA_NS39 + T_N_STRESS;
                when "00101001" => P_EDA_NS40 <= P_EDA_NS40 + T_N_STRESS;
                when "00101010" => P_EDA_NS41 <= P_EDA_NS41 + T_N_STRESS;
                when "00101011" => P_EDA_NS42 <= P_EDA_NS42 + T_N_STRESS;
                when "00101100" => P_EDA_NS43 <= P_EDA_NS43 + T_N_STRESS;
                when "00101101" => P_EDA_NS44 <= P_EDA_NS44 + T_N_STRESS;
                when "00101110" => P_EDA_NS45 <= P_EDA_NS45 + T_N_STRESS;
                when "00101111" => P_EDA_NS46 <= P_EDA_NS46 + T_N_STRESS;
                when "00110000" => P_EDA_NS47 <= P_EDA_NS47 + T_N_STRESS;
                when "00110001" => P_EDA_NS48 <= P_EDA_NS48 + T_N_STRESS;
                when "00110010" => P_EDA_NS49 <= P_EDA_NS49 + T_N_STRESS;
                when "00110011" => P_EDA_NS50 <= P_EDA_NS50 + T_N_STRESS;
                when "00110100" => P_EDA_NS51 <= P_EDA_NS51 + T_N_STRESS;
                when "00110101" => P_EDA_NS52 <= P_EDA_NS52 + T_N_STRESS;
                when "00110110" => P_EDA_NS53 <= P_EDA_NS53 + T_N_STRESS;
                when "00110111" => P_EDA_NS54 <= P_EDA_NS54 + T_N_STRESS;
                when "00111000" => P_EDA_NS55 <= P_EDA_NS55 + T_N_STRESS;
                when "00111001" => P_EDA_NS56 <= P_EDA_NS56 + T_N_STRESS;
                when "00111010" => P_EDA_NS57 <= P_EDA_NS57 + T_N_STRESS;
                when "00111011" => P_EDA_NS58 <= P_EDA_NS58 + T_N_STRESS;
                when "00111100" => P_EDA_NS59 <= P_EDA_NS59 + T_N_STRESS;
                when "00111101" => P_EDA_NS60 <= P_EDA_NS60 + T_N_STRESS;
                when "00111110" => P_EDA_NS61 <= P_EDA_NS61 + T_N_STRESS;
                when "00111111" => P_EDA_NS62 <= P_EDA_NS62 + T_N_STRESS;
                when "01000000" => P_EDA_NS63 <= P_EDA_NS63 + T_N_STRESS;
                when "01000001" => P_EDA_NS64 <= P_EDA_NS64 + T_N_STRESS;
                when "01000010" => P_EDA_NS65 <= P_EDA_NS65 + T_N_STRESS;
                when "01000011" => P_EDA_NS66 <= P_EDA_NS66 + T_N_STRESS;
                when "01000100" => P_EDA_NS67 <= P_EDA_NS67 + T_N_STRESS;
                when "01000101" => P_EDA_NS68 <= P_EDA_NS68 + T_N_STRESS;
                when "01000110" => P_EDA_NS69 <= P_EDA_NS69 + T_N_STRESS;
                when "01000111" => P_EDA_NS70 <= P_EDA_NS70 + T_N_STRESS;
                when "01001000" => P_EDA_NS71 <= P_EDA_NS71 + T_N_STRESS;
                when "01001001" => P_EDA_NS72 <= P_EDA_NS72 + T_N_STRESS;
                when "01001010" => P_EDA_NS73 <= P_EDA_NS73 + T_N_STRESS;
                when "01001011" => P_EDA_NS74 <= P_EDA_NS74 + T_N_STRESS;
                when "01001100" => P_EDA_NS75 <= P_EDA_NS75 + T_N_STRESS;
                when "01001101" => P_EDA_NS76 <= P_EDA_NS76 + T_N_STRESS;
                when "01001110" => P_EDA_NS77 <= P_EDA_NS77 + T_N_STRESS;
                when "01001111" => P_EDA_NS78 <= P_EDA_NS78 + T_N_STRESS;
                when "01010000" => P_EDA_NS79 <= P_EDA_NS79 + T_N_STRESS;
                when "01010001" => P_EDA_NS80 <= P_EDA_NS80 + T_N_STRESS;
                when "01010010" => P_EDA_NS81 <= P_EDA_NS81 + T_N_STRESS;
                when "01010011" => P_EDA_NS82 <= P_EDA_NS82 + T_N_STRESS;
                when "01010100" => P_EDA_NS83 <= P_EDA_NS83 + T_N_STRESS;
                when "01010101" => P_EDA_NS84 <= P_EDA_NS84 + T_N_STRESS;
                when "01010110" => P_EDA_NS85 <= P_EDA_NS85 + T_N_STRESS;
                when "01010111" => P_EDA_NS86 <= P_EDA_NS86 + T_N_STRESS;
                when "01011000" => P_EDA_NS87 <= P_EDA_NS87 + T_N_STRESS;
                when "01011001" => P_EDA_NS88 <= P_EDA_NS88 + T_N_STRESS;
                when "01011010" => P_EDA_NS89 <= P_EDA_NS89 + T_N_STRESS;
                when "01011011" => P_EDA_NS90 <= P_EDA_NS90 + T_N_STRESS;
                when "01011100" => P_EDA_NS91 <= P_EDA_NS91 + T_N_STRESS;
                when "01011101" => P_EDA_NS92 <= P_EDA_NS92 + T_N_STRESS;
                when "01011110" => P_EDA_NS93 <= P_EDA_NS93 + T_N_STRESS;
                when "01011111" => P_EDA_NS94 <= P_EDA_NS94 + T_N_STRESS;
                when "01100000" => P_EDA_NS95 <= P_EDA_NS95 + T_N_STRESS;
                when "01100001" => P_EDA_NS96 <= P_EDA_NS96 + T_N_STRESS;
                when "01100010" => P_EDA_NS97 <= P_EDA_NS97 + T_N_STRESS;
                when "01100011" => P_EDA_NS98 <= P_EDA_NS98 + T_N_STRESS;
                when "01100100" => P_EDA_NS99 <= P_EDA_NS99 + T_N_STRESS;
                when "01100101" => P_EDA_NS100 <= P_EDA_NS100 + T_N_STRESS;
                when "01100110" => P_EDA_NS101 <= P_EDA_NS101 + T_N_STRESS;
                when "01100111" => P_EDA_NS102 <= P_EDA_NS102 + T_N_STRESS;
                when "01101000" => P_EDA_NS103 <= P_EDA_NS103 + T_N_STRESS;
                when "01101001" => P_EDA_NS104 <= P_EDA_NS104 + T_N_STRESS;
                when "01101010" => P_EDA_NS105 <= P_EDA_NS105 + T_N_STRESS;
                when "01101011" => P_EDA_NS106 <= P_EDA_NS106 + T_N_STRESS;
                when "01101100" => P_EDA_NS107 <= P_EDA_NS107 + T_N_STRESS;
                when "10101110" => P_EDA_NS108 <= P_EDA_NS108 + T_N_STRESS;
                when "10101111" => P_EDA_NS109 <= P_EDA_NS109 + T_N_STRESS;
                when "10110000" => P_EDA_NS110 <= P_EDA_NS110 + T_N_STRESS;
				when others            => null;
			end case;
			
		else 
			not_stress_score <= (others => '0');
			P_TEMP_NS <= (others => '0'); 
			P_EDA_NS <= (others => '0');
			P_HR_NS <= (others => '0');
		end if;
	   end if;
	end process;
	


end behavioral;