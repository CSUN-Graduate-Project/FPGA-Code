-----------------------------------------------------------------
-- Created By: Richard Cho
-- Create Date: 3/17/2022
-----------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity SCORE_CALC_T is
    
    port (
        clk : in std_logic; -- system clock
        rst : in std_logic; -- system reset
		temp : in std_logic_vector (8 downto 0); -- celcius
		eda : in std_logic_vector (6 downto 0); --micro siemens
		hr : in std_logic_vector (10 downto 0); -- bpm
		s1 : in std_logic_vector (1 downto 0); -- switch for states
		status : out std_logic_vector (1 downto 0)); -- output
		
end SCORE_CALC_T;

architecture behavioral of SCORE_CALC_T is

	
	
	signal P_TEMP_S1 : unsigned(11 downto 0);
	signal P_TEMP_S2 : unsigned(11 downto 0);
	signal P_TEMP_S3 : unsigned(11 downto 0);
	signal P_TEMP_S4 : unsigned(11 downto 0);
	signal P_TEMP_S5 : unsigned(11 downto 0);
	signal P_TEMP_S6 : unsigned(11 downto 0);
	signal P_TEMP_S7 : unsigned(11 downto 0);
	signal P_TEMP_S8 : unsigned(11 downto 0);
	signal P_TEMP_S9 : unsigned(11 downto 0);
	signal P_TEMP_S10 : unsigned(11 downto 0);
	signal P_TEMP_S11 : unsigned(11 downto 0);
	signal P_TEMP_S12 : unsigned(11 downto 0);
	signal P_TEMP_S13 : unsigned(11 downto 0);
	signal P_TEMP_S14 : unsigned(11 downto 0);
	signal P_TEMP_S15 : unsigned(11 downto 0);
	signal P_TEMP_S16 : unsigned(11 downto 0);
	signal P_TEMP_S17 : unsigned(11 downto 0);
	signal P_TEMP_S18 : unsigned(11 downto 0);
	signal P_TEMP_S19 : unsigned(11 downto 0);
	signal P_TEMP_S20 : unsigned(11 downto 0);
	signal P_TEMP_S21 : unsigned(11 downto 0);
	signal P_TEMP_S22 : unsigned(11 downto 0);
	signal P_TEMP_S23 : unsigned(11 downto 0);
	signal P_TEMP_S24 : unsigned(11 downto 0);
	signal P_TEMP_S25 : unsigned(11 downto 0);
	signal P_TEMP_S26 : unsigned(11 downto 0);
	signal P_TEMP_S27 : unsigned(11 downto 0);
	signal P_TEMP_S28 : unsigned(11 downto 0);
	signal P_TEMP_S29 : unsigned(11 downto 0);
	signal P_TEMP_S30 : unsigned(11 downto 0);
	
	signal P_EDA_S1 : unsigned(11 downto 0);
	signal P_EDA_S2 : unsigned(11 downto 0);
	signal P_EDA_S3 : unsigned(11 downto 0);
	signal P_EDA_S4 : unsigned(11 downto 0);
	signal P_EDA_S5 : unsigned(11 downto 0);
	signal P_EDA_S6 : unsigned(11 downto 0);
	signal P_EDA_S7 : unsigned(11 downto 0);
	signal P_EDA_S8 : unsigned(11 downto 0);
	signal P_EDA_S9 : unsigned(11 downto 0);
	signal P_EDA_S10 : unsigned(11 downto 0);
	signal P_EDA_S11 : unsigned(11 downto 0);
	signal P_EDA_S12 : unsigned(11 downto 0);
	signal P_EDA_S13 : unsigned(11 downto 0);
	signal P_EDA_S14 : unsigned(11 downto 0);
	signal P_EDA_S15 : unsigned(11 downto 0);
	signal P_EDA_S16 : unsigned(11 downto 0);
	signal P_EDA_S17 : unsigned(11 downto 0);
	signal P_EDA_S18 : unsigned(11 downto 0);
	signal P_EDA_S19 : unsigned(11 downto 0);
	signal P_EDA_S20 : unsigned(11 downto 0);
	signal P_EDA_S21 : unsigned(11 downto 0);
	signal P_EDA_S22 : unsigned(11 downto 0);
	signal P_EDA_S23 : unsigned(11 downto 0);
	signal P_EDA_S24 : unsigned(11 downto 0);
	signal P_EDA_S25 : unsigned(11 downto 0);
	signal P_EDA_S26 : unsigned(11 downto 0);
	signal P_EDA_S27 : unsigned(11 downto 0);
	signal P_EDA_S28 : unsigned(11 downto 0);
	signal P_EDA_S29 : unsigned(11 downto 0);
	signal P_EDA_S30 : unsigned(11 downto 0);
	signal P_EDA_S31 : unsigned(11 downto 0);
	signal P_EDA_S32 : unsigned(11 downto 0);
	signal P_EDA_S33 : unsigned(11 downto 0);
	signal P_EDA_S34 : unsigned(11 downto 0);
	signal P_EDA_S35 : unsigned(11 downto 0);
	signal P_EDA_S36 : unsigned(11 downto 0);
	signal P_EDA_S37 : unsigned(11 downto 0);
	signal P_EDA_S38 : unsigned(11 downto 0);
	signal P_EDA_S39 : unsigned(11 downto 0);
	signal P_EDA_S40 : unsigned(11 downto 0);
	signal P_EDA_S41 : unsigned(11 downto 0);
	signal P_EDA_S42 : unsigned(11 downto 0);
	signal P_EDA_S43 : unsigned(11 downto 0);
	signal P_EDA_S44 : unsigned(11 downto 0);
	signal P_EDA_S45 : unsigned(11 downto 0);
	signal P_EDA_S46 : unsigned(11 downto 0);
	signal P_EDA_S47 : unsigned(11 downto 0);
	signal P_EDA_S48 : unsigned(11 downto 0);
	signal P_EDA_S49 : unsigned(11 downto 0);
	signal P_EDA_S50 : unsigned(11 downto 0);
	signal P_EDA_S51 : unsigned(11 downto 0);
	signal P_EDA_S52 : unsigned(11 downto 0);
	signal P_EDA_S53 : unsigned(11 downto 0);
	signal P_EDA_S54 : unsigned(11 downto 0);
	signal P_EDA_S55 : unsigned(11 downto 0);
	signal P_EDA_S56 : unsigned(11 downto 0);
	signal P_EDA_S57 : unsigned(11 downto 0);
	signal P_EDA_S58 : unsigned(11 downto 0);
	signal P_EDA_S59 : unsigned(11 downto 0);
	signal P_EDA_S60 : unsigned(11 downto 0);
	signal P_EDA_S61 : unsigned(11 downto 0);
	signal P_EDA_S62 : unsigned(11 downto 0);
	signal P_EDA_S63 : unsigned(11 downto 0);
	signal P_EDA_S64 : unsigned(11 downto 0);
	signal P_EDA_S65 : unsigned(11 downto 0);
	
	
	signal P_HR_S1 : unsigned(11 downto 0); 
	signal P_HR_S2 : unsigned(11 downto 0); 
	signal P_HR_S3 : unsigned(11 downto 0); 
	signal P_HR_S4 : unsigned(11 downto 0); 
	signal P_HR_S5 : unsigned(11 downto 0); 
	signal P_HR_S6 : unsigned(11 downto 0); 
	signal P_HR_S7 : unsigned(11 downto 0); 
	signal P_HR_S8 : unsigned(11 downto 0); 
	signal P_HR_S9 : unsigned(11 downto 0); 
	signal P_HR_S10 : unsigned(11 downto 0);
	signal P_HR_S11 : unsigned(11 downto 0);
	signal P_HR_S12 : unsigned(11 downto 0);
	signal P_HR_S13 : unsigned(11 downto 0);
	signal P_HR_S14 : unsigned(11 downto 0);
	signal P_HR_S15 : unsigned(11 downto 0);
	signal P_HR_S16 : unsigned(11 downto 0);
	signal P_HR_S17 : unsigned(11 downto 0);
	signal P_HR_S18 : unsigned(11 downto 0);
	signal P_HR_S19 : unsigned(11 downto 0);
	signal P_HR_S20 : unsigned(11 downto 0);
	signal P_HR_S21 : unsigned(11 downto 0);
	signal P_HR_S22 : unsigned(11 downto 0);
	signal P_HR_S23 : unsigned(11 downto 0);
	signal P_HR_S24 : unsigned(11 downto 0);
	signal P_HR_S25 : unsigned(11 downto 0);
	signal P_HR_S26 : unsigned(11 downto 0);
	signal P_HR_S27 : unsigned(11 downto 0);
	signal P_HR_S28 : unsigned(11 downto 0);
	signal P_HR_S29 : unsigned(11 downto 0);
	signal P_HR_S30 : unsigned(11 downto 0);
	signal P_HR_S31 : unsigned(11 downto 0);
	signal P_HR_S32 : unsigned(11 downto 0);
	signal P_HR_S33 : unsigned(11 downto 0);
	signal P_HR_S34 : unsigned(11 downto 0);
	signal P_HR_S35 : unsigned(11 downto 0);
	signal P_HR_S36 : unsigned(11 downto 0);
	signal P_HR_S37 : unsigned(11 downto 0);
	signal P_HR_S38 : unsigned(11 downto 0);
	signal P_HR_S39 : unsigned(11 downto 0);
	signal P_HR_S40 : unsigned(11 downto 0);
	signal P_HR_S41 : unsigned(11 downto 0);
	signal P_HR_S42 : unsigned(11 downto 0);
	signal P_HR_S43 : unsigned(11 downto 0);
	signal P_HR_S44 : unsigned(11 downto 0);
	signal P_HR_S45 : unsigned(11 downto 0);
	signal P_HR_S46 : unsigned(11 downto 0);
	signal P_HR_S47 : unsigned(11 downto 0);
	signal P_HR_S48 : unsigned(11 downto 0);
	signal P_HR_S49 : unsigned(11 downto 0);
	signal P_HR_S50 : unsigned(11 downto 0);
	signal P_HR_S51 : unsigned(11 downto 0);
	signal P_HR_S52 : unsigned(11 downto 0);
	signal P_HR_S53 : unsigned(11 downto 0);
	signal P_HR_S54 : unsigned(11 downto 0);
	signal P_HR_S55 : unsigned(11 downto 0);
	signal P_HR_S56 : unsigned(11 downto 0);
	signal P_HR_S57 : unsigned(11 downto 0);
	signal P_HR_S58 : unsigned(11 downto 0);
	signal P_HR_S59 : unsigned(11 downto 0);
	signal P_HR_S60 : unsigned(11 downto 0);
	signal P_HR_S61 : unsigned(11 downto 0);
	signal P_HR_S62 : unsigned(11 downto 0);
	signal P_HR_S63 : unsigned(11 downto 0);
	signal P_HR_S64 : unsigned(11 downto 0);
	signal P_HR_S65 : unsigned(11 downto 0);
	signal P_HR_S66 : unsigned(11 downto 0);
	signal P_HR_S67 : unsigned(11 downto 0);
	signal P_HR_S68 : unsigned(11 downto 0);
	signal P_HR_S69 : unsigned(11 downto 0);
	signal P_HR_S70 : unsigned(11 downto 0);
	signal P_HR_S71 : unsigned(11 downto 0);
	signal P_HR_S72 : unsigned(11 downto 0);
	signal P_HR_S73 : unsigned(11 downto 0);
	signal P_HR_S74 : unsigned(11 downto 0);
	signal P_HR_S75 : unsigned(11 downto 0);
	signal P_HR_S76 : unsigned(11 downto 0);
	signal P_HR_S77 : unsigned(11 downto 0);
	signal P_HR_S78 : unsigned(11 downto 0);
	signal P_HR_S79 : unsigned(11 downto 0);
	signal P_HR_S80 : unsigned(11 downto 0);
	signal P_HR_S81 : unsigned(11 downto 0);
	signal P_HR_S82 : unsigned(11 downto 0);
	signal P_HR_S83 : unsigned(11 downto 0);
	signal P_HR_S84 : unsigned(11 downto 0);
	signal P_HR_S85 : unsigned(11 downto 0);
	signal P_HR_S86 : unsigned(11 downto 0);
	signal P_HR_S87 : unsigned(11 downto 0);
	signal P_HR_S88 : unsigned(11 downto 0);
	signal P_HR_S89 : unsigned(11 downto 0);
	signal P_HR_S90 : unsigned(11 downto 0);
	signal P_HR_S91 : unsigned(11 downto 0);
	signal P_HR_S92 : unsigned(11 downto 0);
	signal P_HR_S93 : unsigned(11 downto 0);
	signal P_HR_S94 : unsigned(11 downto 0);
	signal P_HR_S95 : unsigned(11 downto 0);
	signal P_HR_S96 : unsigned(11 downto 0);
	signal P_HR_S97 : unsigned(11 downto 0);
	signal P_HR_S98 : unsigned(11 downto 0);
	signal P_HR_S99 : unsigned(11 downto 0);
	signal P_HR_S100 : unsigned(11 downto 0);
	signal P_HR_S101 : unsigned(11 downto 0);
	signal P_HR_S102 : unsigned(11 downto 0);
	signal P_HR_S103 : unsigned(11 downto 0);
	signal P_HR_S104 : unsigned(11 downto 0);
	signal P_HR_S105 : unsigned(11 downto 0);
	signal P_HR_S106 : unsigned(11 downto 0);
	signal P_HR_S107 : unsigned(11 downto 0);
	signal P_HR_S108 : unsigned(11 downto 0);
	signal P_HR_S109 : unsigned(11 downto 0);
	signal P_HR_S110 : unsigned(11 downto 0);
	signal P_HR_S111 : unsigned(11 downto 0);
	signal P_HR_S112 : unsigned(11 downto 0);
	signal P_HR_S113 : unsigned(11 downto 0);
	signal P_HR_S114 : unsigned(11 downto 0);
	signal P_HR_S115 : unsigned(11 downto 0);
	signal P_HR_S116 : unsigned(11 downto 0);
	signal P_HR_S117 : unsigned(11 downto 0);
	signal P_HR_S118 : unsigned(11 downto 0);
	signal P_HR_S119 : unsigned(11 downto 0);
	signal P_HR_S120 : unsigned(11 downto 0);
	signal P_HR_S121 : unsigned(11 downto 0);
	signal P_HR_S122 : unsigned(11 downto 0);
	signal P_HR_S123 : unsigned(11 downto 0);
	signal P_HR_S124 : unsigned(11 downto 0);
	signal P_HR_S125 : unsigned(11 downto 0);
	signal P_HR_S126 : unsigned(11 downto 0);
	signal P_HR_S127 : unsigned(11 downto 0);
	signal P_HR_S128 : unsigned(11 downto 0);
	signal P_HR_S129 : unsigned(11 downto 0);
	signal P_HR_S130 : unsigned(11 downto 0);
	signal P_HR_S131 : unsigned(11 downto 0);
	signal P_HR_S132 : unsigned(11 downto 0);
	signal P_HR_S133 : unsigned(11 downto 0);
	signal P_HR_S134 : unsigned(11 downto 0);
	signal P_HR_S135 : unsigned(11 downto 0);
	signal P_HR_S136 : unsigned(11 downto 0);
	signal P_HR_S137 : unsigned(11 downto 0);
	signal P_HR_S138 : unsigned(11 downto 0);
	signal P_HR_S139 : unsigned(11 downto 0);
	signal P_HR_S140 : unsigned(11 downto 0);
	signal P_HR_S141 : unsigned(11 downto 0);
	signal P_HR_S142 : unsigned(11 downto 0);
	signal P_HR_S143 : unsigned(11 downto 0);
	signal P_HR_S144 : unsigned(11 downto 0);
	signal P_HR_S145 : unsigned(11 downto 0);
	signal P_HR_S146 : unsigned(11 downto 0);
	signal P_HR_S147 : unsigned(11 downto 0);
	signal P_HR_S148 : unsigned(11 downto 0);
	signal P_HR_S149 : unsigned(11 downto 0);
	signal P_HR_S150 : unsigned(11 downto 0);
	signal P_HR_S151 : unsigned(11 downto 0);
	signal P_HR_S152 : unsigned(11 downto 0);
	signal P_HR_S153 : unsigned(11 downto 0);
	signal P_HR_S154 : unsigned(11 downto 0);
	signal P_HR_S155 : unsigned(11 downto 0);
	signal P_HR_S156 : unsigned(11 downto 0);
	signal P_HR_S157 : unsigned(11 downto 0);
	signal P_HR_S158 : unsigned(11 downto 0);
	signal P_HR_S159 : unsigned(11 downto 0);
	signal P_HR_S160 : unsigned(11 downto 0);
	signal P_HR_S161 : unsigned(11 downto 0);
	signal P_HR_S162 : unsigned(11 downto 0);
	signal P_HR_S163 : unsigned(11 downto 0);
	signal P_HR_S164 : unsigned(11 downto 0);
	signal P_HR_S165 : unsigned(11 downto 0);
	signal P_HR_S166 : unsigned(11 downto 0);
	signal P_HR_S167 : unsigned(11 downto 0);
	signal P_HR_S168 : unsigned(11 downto 0);
	signal P_HR_S169 : unsigned(11 downto 0);
	signal P_HR_S170 : unsigned(11 downto 0);
	signal P_HR_S171 : unsigned(11 downto 0);
	signal P_HR_S172 : unsigned(11 downto 0);
	signal P_HR_S173 : unsigned(11 downto 0);
	signal P_HR_S174 : unsigned(11 downto 0);
	signal P_HR_S175 : unsigned(11 downto 0);
	signal P_HR_S176 : unsigned(11 downto 0);
	signal P_HR_S177 : unsigned(11 downto 0);
	signal P_HR_S178 : unsigned(11 downto 0);
	signal P_HR_S179 : unsigned(11 downto 0);
	signal P_HR_S180 : unsigned(11 downto 0);
	signal P_HR_S181 : unsigned(11 downto 0);
	signal P_HR_S182 : unsigned(11 downto 0);
	signal P_HR_S183 : unsigned(11 downto 0);
	signal P_HR_S184 : unsigned(11 downto 0);
	signal P_HR_S185 : unsigned(11 downto 0);
	signal P_HR_S186 : unsigned(11 downto 0);
	signal P_HR_S187 : unsigned(11 downto 0);
	signal P_HR_S188 : unsigned(11 downto 0);
	signal P_HR_S189 : unsigned(11 downto 0);
	signal P_HR_S190 : unsigned(11 downto 0);
	signal P_HR_S191 : unsigned(11 downto 0);
	signal P_HR_S192 : unsigned(11 downto 0);
	signal P_HR_S193 : unsigned(11 downto 0);
	signal P_HR_S194 : unsigned(11 downto 0);
	signal P_HR_S195 : unsigned(11 downto 0);
	signal P_HR_S196 : unsigned(11 downto 0);
	signal P_HR_S197 : unsigned(11 downto 0);
	signal P_HR_S198 : unsigned(11 downto 0);
	signal P_HR_S199 : unsigned(11 downto 0);
	signal P_HR_S200 : unsigned(11 downto 0);
	signal P_HR_S201 : unsigned(11 downto 0);
	signal P_HR_S202 : unsigned(11 downto 0);
	signal P_HR_S203 : unsigned(11 downto 0);
	signal P_HR_S204 : unsigned(11 downto 0);
	signal P_HR_S205 : unsigned(11 downto 0);
	signal P_HR_S206 : unsigned(11 downto 0);
	signal P_HR_S207 : unsigned(11 downto 0);
	signal P_HR_S208 : unsigned(11 downto 0);
	signal P_HR_S209 : unsigned(11 downto 0);
	signal P_HR_S210 : unsigned(11 downto 0);
	signal P_HR_S211 : unsigned(11 downto 0);
	signal P_HR_S212 : unsigned(11 downto 0);
	signal P_HR_S213 : unsigned(11 downto 0);
	signal P_HR_S214 : unsigned(11 downto 0);
	signal P_HR_S215 : unsigned(11 downto 0);
	signal P_HR_S216 : unsigned(11 downto 0);
	signal P_HR_S217 : unsigned(11 downto 0);
	signal P_HR_S218 : unsigned(11 downto 0);
	signal P_HR_S219 : unsigned(11 downto 0);
	signal P_HR_S220 : unsigned(11 downto 0);
	signal P_HR_S221 : unsigned(11 downto 0);
	signal P_HR_S222 : unsigned(11 downto 0);
	signal P_HR_S223 : unsigned(11 downto 0);
	signal P_HR_S224 : unsigned(11 downto 0);
	signal P_HR_S225 : unsigned(11 downto 0);
	signal P_HR_S226 : unsigned(11 downto 0);
	signal P_HR_S227 : unsigned(11 downto 0);
	signal P_HR_S228 : unsigned(11 downto 0);
	signal P_HR_S229 : unsigned(11 downto 0);
	signal P_HR_S230 : unsigned(11 downto 0);
	signal P_HR_S231 : unsigned(11 downto 0);
	signal P_HR_S232 : unsigned(11 downto 0);
	signal P_HR_S233 : unsigned(11 downto 0);
	signal P_HR_S234 : unsigned(11 downto 0);
	signal P_HR_S235 : unsigned(11 downto 0);
	signal P_HR_S236 : unsigned(11 downto 0);
	signal P_HR_S237 : unsigned(11 downto 0);
	signal P_HR_S238 : unsigned(11 downto 0);
	signal P_HR_S239 : unsigned(11 downto 0);
	signal P_HR_S240 : unsigned(11 downto 0);
	signal P_HR_S241 : unsigned(11 downto 0);
	signal P_HR_S242 : unsigned(11 downto 0);
	signal P_HR_S243 : unsigned(11 downto 0);
	signal P_HR_S244 : unsigned(11 downto 0);
	signal P_HR_S245 : unsigned(11 downto 0);
	signal P_HR_S246 : unsigned(11 downto 0);
	signal P_HR_S247 : unsigned(11 downto 0);
	signal P_HR_S248 : unsigned(11 downto 0);
	signal P_HR_S249 : unsigned(11 downto 0);
	signal P_HR_S250 : unsigned(11 downto 0);
	signal P_HR_S251 : unsigned(11 downto 0);
	signal P_HR_S252 : unsigned(11 downto 0);
	signal P_HR_S253 : unsigned(11 downto 0);
	signal P_HR_S254 : unsigned(11 downto 0);
	signal P_HR_S255 : unsigned(11 downto 0);
	signal P_HR_S256 : unsigned(11 downto 0);
	signal P_HR_S257 : unsigned(11 downto 0);
	signal P_HR_S258 : unsigned(11 downto 0);
	signal P_HR_S259 : unsigned(11 downto 0);
	signal P_HR_S260 : unsigned(11 downto 0);
	signal P_HR_S261 : unsigned(11 downto 0);
	signal P_HR_S262 : unsigned(11 downto 0);
	signal P_HR_S263 : unsigned(11 downto 0);
	signal P_HR_S264 : unsigned(11 downto 0);
	signal P_HR_S265 : unsigned(11 downto 0);
	signal P_HR_S266 : unsigned(11 downto 0);
	signal P_HR_S267 : unsigned(11 downto 0);
	signal P_HR_S268 : unsigned(11 downto 0);
	signal P_HR_S269 : unsigned(11 downto 0);
	signal P_HR_S270 : unsigned(11 downto 0);
	signal P_HR_S271 : unsigned(11 downto 0);
	signal P_HR_S272 : unsigned(11 downto 0);
	signal P_HR_S273 : unsigned(11 downto 0);
	signal P_HR_S274 : unsigned(11 downto 0);
	signal P_HR_S275 : unsigned(11 downto 0);
	signal P_HR_S276 : unsigned(11 downto 0);
	signal P_HR_S277 : unsigned(11 downto 0);
	signal P_HR_S278 : unsigned(11 downto 0);
	signal P_HR_S279 : unsigned(11 downto 0);
	signal P_HR_S280 : unsigned(11 downto 0);
	signal P_HR_S281 : unsigned(11 downto 0);
	signal P_HR_S282 : unsigned(11 downto 0);
	signal P_HR_S283 : unsigned(11 downto 0);
	signal P_HR_S284 : unsigned(11 downto 0);
	signal P_HR_S285 : unsigned(11 downto 0);
	signal P_HR_S286 : unsigned(11 downto 0);
	signal P_HR_S287 : unsigned(11 downto 0);
	signal P_HR_S288 : unsigned(11 downto 0);
	signal P_HR_S289 : unsigned(11 downto 0);
	signal P_HR_S290 : unsigned(11 downto 0);
	signal P_HR_S291 : unsigned(11 downto 0);
	signal P_HR_S292 : unsigned(11 downto 0);
	signal P_HR_S293 : unsigned(11 downto 0);
	signal P_HR_S294 : unsigned(11 downto 0);
	signal P_HR_S295 : unsigned(11 downto 0);
	signal P_HR_S296 : unsigned(11 downto 0);
	signal P_HR_S297 : unsigned(11 downto 0);
	signal P_HR_S298 : unsigned(11 downto 0);
	signal P_HR_S299 : unsigned(11 downto 0);
	signal P_HR_S300 : unsigned(11 downto 0);
	signal P_HR_S301 : unsigned(11 downto 0);
	signal P_HR_S302 : unsigned(11 downto 0);
	signal P_HR_S303 : unsigned(11 downto 0);
	signal P_HR_S304 : unsigned(11 downto 0);
	signal P_HR_S305 : unsigned(11 downto 0);
	signal P_HR_S306 : unsigned(11 downto 0);
	signal P_HR_S307 : unsigned(11 downto 0);
	signal P_HR_S308 : unsigned(11 downto 0);
	signal P_HR_S309 : unsigned(11 downto 0);
	signal P_HR_S310 : unsigned(11 downto 0);
	signal P_HR_S311 : unsigned(11 downto 0);
	signal P_HR_S312 : unsigned(11 downto 0);
	signal P_HR_S313 : unsigned(11 downto 0);
	signal P_HR_S314 : unsigned(11 downto 0);
	signal P_HR_S315 : unsigned(11 downto 0);
	signal P_HR_S316 : unsigned(11 downto 0);
	signal P_HR_S317 : unsigned(11 downto 0);
	signal P_HR_S318 : unsigned(11 downto 0);
	signal P_HR_S319 : unsigned(11 downto 0);
	signal P_HR_S320 : unsigned(11 downto 0);
	signal P_HR_S321 : unsigned(11 downto 0);
	signal P_HR_S322 : unsigned(11 downto 0);
	signal P_HR_S323 : unsigned(11 downto 0);
	signal P_HR_S324 : unsigned(11 downto 0);
	signal P_HR_S325 : unsigned(11 downto 0);
	signal P_HR_S326 : unsigned(11 downto 0);
	signal P_HR_S327 : unsigned(11 downto 0);
	signal P_HR_S328 : unsigned(11 downto 0);
	signal P_HR_S329 : unsigned(11 downto 0);
	signal P_HR_S330 : unsigned(11 downto 0);
	signal P_HR_S331 : unsigned(11 downto 0);
	signal P_HR_S332 : unsigned(11 downto 0);
	signal P_HR_S333 : unsigned(11 downto 0);
	signal P_HR_S334 : unsigned(11 downto 0);
	signal P_HR_S335 : unsigned(11 downto 0);
	signal P_HR_S336 : unsigned(11 downto 0);
	signal P_HR_S337 : unsigned(11 downto 0);
	signal P_HR_S338 : unsigned(11 downto 0);
	signal P_HR_S339 : unsigned(11 downto 0);
	signal P_HR_S340 : unsigned(11 downto 0);
	signal P_HR_S341 : unsigned(11 downto 0);
	signal P_HR_S342 : unsigned(11 downto 0);
	signal P_HR_S343 : unsigned(11 downto 0);
	signal P_HR_S344 : unsigned(11 downto 0);
	signal P_HR_S345 : unsigned(11 downto 0);
	signal P_HR_S346 : unsigned(11 downto 0);
	signal P_HR_S347 : unsigned(11 downto 0);
	signal P_HR_S348 : unsigned(11 downto 0);
	signal P_HR_S349 : unsigned(11 downto 0);
	signal P_HR_S350 : unsigned(11 downto 0);
	signal P_HR_S351 : unsigned(11 downto 0);
	signal P_HR_S352 : unsigned(11 downto 0);
	signal P_HR_S353 : unsigned(11 downto 0);
	signal P_HR_S354 : unsigned(11 downto 0);
	signal P_HR_S355 : unsigned(11 downto 0);
	signal P_HR_S356 : unsigned(11 downto 0);
	signal P_HR_S357 : unsigned(11 downto 0);
	signal P_HR_S358 : unsigned(11 downto 0);
	signal P_HR_S359 : unsigned(11 downto 0);
	signal P_HR_S360 : unsigned(11 downto 0);
	signal P_HR_S361 : unsigned(11 downto 0);
	signal P_HR_S362 : unsigned(11 downto 0);
	signal P_HR_S363 : unsigned(11 downto 0);
	signal P_HR_S364 : unsigned(11 downto 0);
	signal P_HR_S365 : unsigned(11 downto 0);
	signal P_HR_S366 : unsigned(11 downto 0);
	signal P_HR_S367 : unsigned(11 downto 0);
	signal P_HR_S368 : unsigned(11 downto 0);
	signal P_HR_S369 : unsigned(11 downto 0);
	signal P_HR_S370 : unsigned(11 downto 0);
	signal P_HR_S371 : unsigned(11 downto 0);
	signal P_HR_S372 : unsigned(11 downto 0);
	signal P_HR_S373 : unsigned(11 downto 0);
	signal P_HR_S374 : unsigned(11 downto 0);
	signal P_HR_S375 : unsigned(11 downto 0);
	signal P_HR_S376 : unsigned(11 downto 0);
	signal P_HR_S377 : unsigned(11 downto 0);
	signal P_HR_S378 : unsigned(11 downto 0);
	signal P_HR_S379 : unsigned(11 downto 0);
	signal P_HR_S380 : unsigned(11 downto 0);
	signal P_HR_S381 : unsigned(11 downto 0);
	signal P_HR_S382 : unsigned(11 downto 0);
	signal P_HR_S383 : unsigned(11 downto 0);
	signal P_HR_S384 : unsigned(11 downto 0);
	signal P_HR_S385 : unsigned(11 downto 0);
	signal P_HR_S386 : unsigned(11 downto 0);
	signal P_HR_S387 : unsigned(11 downto 0);
	signal P_HR_S388 : unsigned(11 downto 0);
	signal P_HR_S389 : unsigned(11 downto 0);
	signal P_HR_S390 : unsigned(11 downto 0);
	signal P_HR_S391 : unsigned(11 downto 0);
	signal P_HR_S392 : unsigned(11 downto 0);
	signal P_HR_S393 : unsigned(11 downto 0);
	signal P_HR_S394 : unsigned(11 downto 0);
	signal P_HR_S395 : unsigned(11 downto 0);
	signal P_HR_S396 : unsigned(11 downto 0);
	signal P_HR_S397 : unsigned(11 downto 0);
	signal P_HR_S398 : unsigned(11 downto 0);
	signal P_HR_S399 : unsigned(11 downto 0);
	signal P_HR_S400 : unsigned(11 downto 0);
	signal P_HR_S401 : unsigned(11 downto 0);
	signal P_HR_S402 : unsigned(11 downto 0);
	signal P_HR_S403 : unsigned(11 downto 0);
	signal P_HR_S404 : unsigned(11 downto 0);
	signal P_HR_S405 : unsigned(11 downto 0);
	signal P_HR_S406 : unsigned(11 downto 0);
	signal P_HR_S407 : unsigned(11 downto 0);
	signal P_HR_S408 : unsigned(11 downto 0);
	signal P_HR_S409 : unsigned(11 downto 0);
	signal P_HR_S410 : unsigned(11 downto 0);
	signal P_HR_S411 : unsigned(11 downto 0);
	signal P_HR_S412 : unsigned(11 downto 0);
	signal P_HR_S413 : unsigned(11 downto 0);
	signal P_HR_S414 : unsigned(11 downto 0);
	signal P_HR_S415 : unsigned(11 downto 0);
	signal P_HR_S416 : unsigned(11 downto 0);
	signal P_HR_S417 : unsigned(11 downto 0);
	signal P_HR_S418 : unsigned(11 downto 0);
	signal P_HR_S419 : unsigned(11 downto 0);
	signal P_HR_S420 : unsigned(11 downto 0);
	signal P_HR_S421 : unsigned(11 downto 0);
	signal P_HR_S422 : unsigned(11 downto 0);
	signal P_HR_S423 : unsigned(11 downto 0);
	signal P_HR_S424 : unsigned(11 downto 0);
	signal P_HR_S425 : unsigned(11 downto 0);
	signal P_HR_S426 : unsigned(11 downto 0);
	signal P_HR_S427 : unsigned(11 downto 0);
	signal P_HR_S428 : unsigned(11 downto 0);
	
	signal P_TEMP_NS1 : unsigned(11 downto 0);
	signal P_TEMP_NS2 : unsigned(11 downto 0);
	signal P_TEMP_NS3 : unsigned(11 downto 0);
	signal P_TEMP_NS4 : unsigned(11 downto 0);
	signal P_TEMP_NS5 : unsigned(11 downto 0);
	signal P_TEMP_NS6 : unsigned(11 downto 0);
	signal P_TEMP_NS7 : unsigned(11 downto 0);
	signal P_TEMP_NS8 : unsigned(11 downto 0);
	signal P_TEMP_NS9 : unsigned(11 downto 0);
	signal P_TEMP_NS10 : unsigned(11 downto 0);
	signal P_TEMP_NS11 : unsigned(11 downto 0);
	signal P_TEMP_NS12 : unsigned(11 downto 0);
	signal P_TEMP_NS13 : unsigned(11 downto 0);
	signal P_TEMP_NS14 : unsigned(11 downto 0);
	signal P_TEMP_NS15 : unsigned(11 downto 0);
	signal P_TEMP_NS16 : unsigned(11 downto 0);
	signal P_TEMP_NS17 : unsigned(11 downto 0);
	signal P_TEMP_NS18 : unsigned(11 downto 0);
	signal P_TEMP_NS19 : unsigned(11 downto 0);
	signal P_TEMP_NS20 : unsigned(11 downto 0);
	signal P_TEMP_NS21 : unsigned(11 downto 0);
	signal P_TEMP_NS22 : unsigned(11 downto 0);
	signal P_TEMP_NS23 : unsigned(11 downto 0);
	signal P_TEMP_NS24 : unsigned(11 downto 0);
	signal P_TEMP_NS25 : unsigned(11 downto 0);
	signal P_TEMP_NS26 : unsigned(11 downto 0);
	signal P_TEMP_NS27 : unsigned(11 downto 0);
	signal P_TEMP_NS28 : unsigned(11 downto 0);
	signal P_TEMP_NS29 : unsigned(11 downto 0);
	signal P_TEMP_NS30 : unsigned(11 downto 0);
	signal P_TEMP_NS31 : unsigned(11 downto 0);
	signal P_TEMP_NS32 : unsigned(11 downto 0);
	signal P_TEMP_NS33 : unsigned(11 downto 0);
	signal P_TEMP_NS34 : unsigned(11 downto 0);
	signal P_TEMP_NS35 : unsigned(11 downto 0);
	signal P_TEMP_NS36 : unsigned(11 downto 0);
	signal P_TEMP_NS37 : unsigned(11 downto 0);
	signal P_TEMP_NS38 : unsigned(11 downto 0);
	signal P_TEMP_NS39 : unsigned(11 downto 0);
	signal P_TEMP_NS40 : unsigned(11 downto 0);
	signal P_TEMP_NS41 : unsigned(11 downto 0);
	signal P_TEMP_NS42 : unsigned(11 downto 0);
	signal P_TEMP_NS43 : unsigned(11 downto 0);
	signal P_TEMP_NS44 : unsigned(11 downto 0);
	signal P_TEMP_NS45 : unsigned(11 downto 0);
	signal P_TEMP_NS46 : unsigned(11 downto 0);
	signal P_TEMP_NS47 : unsigned(11 downto 0);
	signal P_TEMP_NS48 : unsigned(11 downto 0);
	signal P_TEMP_NS49 : unsigned(11 downto 0);
	signal P_TEMP_NS50 : unsigned(11 downto 0);
	signal P_TEMP_NS51 : unsigned(11 downto 0);
	signal P_TEMP_NS52 : unsigned(11 downto 0);
		
	signal P_HR_NS1 : unsigned(11 downto 0);
	signal P_HR_NS2 : unsigned(11 downto 0);
	signal P_HR_NS3 : unsigned(11 downto 0);
	signal P_HR_NS4 : unsigned(11 downto 0);
	signal P_HR_NS5 : unsigned(11 downto 0);
	signal P_HR_NS6 : unsigned(11 downto 0);
	signal P_HR_NS7 : unsigned(11 downto 0);
	signal P_HR_NS8 : unsigned(11 downto 0);
	signal P_HR_NS9 : unsigned(11 downto 0);
	signal P_HR_NS10 : unsigned(11 downto 0);
	signal P_HR_NS11 : unsigned(11 downto 0);
	signal P_HR_NS12 : unsigned(11 downto 0);
	signal P_HR_NS13 : unsigned(11 downto 0);
	signal P_HR_NS14 : unsigned(11 downto 0);
	signal P_HR_NS15 : unsigned(11 downto 0);
	signal P_HR_NS16 : unsigned(11 downto 0);
	signal P_HR_NS17 : unsigned(11 downto 0);
	signal P_HR_NS18 : unsigned(11 downto 0);
	signal P_HR_NS19 : unsigned(11 downto 0);
	signal P_HR_NS20 : unsigned(11 downto 0);
	signal P_HR_NS21 : unsigned(11 downto 0);
	signal P_HR_NS22 : unsigned(11 downto 0);
	signal P_HR_NS23 : unsigned(11 downto 0);
	signal P_HR_NS24 : unsigned(11 downto 0);
	signal P_HR_NS25 : unsigned(11 downto 0);
	signal P_HR_NS26 : unsigned(11 downto 0);
	signal P_HR_NS27 : unsigned(11 downto 0);
	signal P_HR_NS28 : unsigned(11 downto 0);
	signal P_HR_NS29 : unsigned(11 downto 0);
	signal P_HR_NS30 : unsigned(11 downto 0);
	signal P_HR_NS31 : unsigned(11 downto 0);
	signal P_HR_NS32 : unsigned(11 downto 0);
	signal P_HR_NS33 : unsigned(11 downto 0);
	signal P_HR_NS34 : unsigned(11 downto 0);
	signal P_HR_NS35 : unsigned(11 downto 0);
	signal P_HR_NS36 : unsigned(11 downto 0);
	signal P_HR_NS37 : unsigned(11 downto 0);
	signal P_HR_NS38 : unsigned(11 downto 0);
	signal P_HR_NS39 : unsigned(11 downto 0);
	signal P_HR_NS40 : unsigned(11 downto 0);
	signal P_HR_NS41 : unsigned(11 downto 0);
	signal P_HR_NS42 : unsigned(11 downto 0);
	signal P_HR_NS43 : unsigned(11 downto 0);
	signal P_HR_NS44 : unsigned(11 downto 0);
	signal P_HR_NS45 : unsigned(11 downto 0);
	signal P_HR_NS46 : unsigned(11 downto 0);
	signal P_HR_NS47 : unsigned(11 downto 0);
	signal P_HR_NS48 : unsigned(11 downto 0);
	signal P_HR_NS49 : unsigned(11 downto 0);
	signal P_HR_NS50 : unsigned(11 downto 0);
	signal P_HR_NS51 : unsigned(11 downto 0);
	signal P_HR_NS52 : unsigned(11 downto 0);
	signal P_HR_NS53 : unsigned(11 downto 0);
	signal P_HR_NS54 : unsigned(11 downto 0);
	signal P_HR_NS55 : unsigned(11 downto 0);
	signal P_HR_NS56 : unsigned(11 downto 0);
	signal P_HR_NS57 : unsigned(11 downto 0);
	signal P_HR_NS58 : unsigned(11 downto 0);
	signal P_HR_NS59 : unsigned(11 downto 0);
	signal P_HR_NS60 : unsigned(11 downto 0);
	signal P_HR_NS61 : unsigned(11 downto 0);
	signal P_HR_NS62 : unsigned(11 downto 0);
	signal P_HR_NS63 : unsigned(11 downto 0);
	signal P_HR_NS64 : unsigned(11 downto 0);
	signal P_HR_NS65 : unsigned(11 downto 0);
	signal P_HR_NS66 : unsigned(11 downto 0);
	signal P_HR_NS67 : unsigned(11 downto 0);
	signal P_HR_NS68 : unsigned(11 downto 0);
	signal P_HR_NS69 : unsigned(11 downto 0);
	signal P_HR_NS70 : unsigned(11 downto 0);
	signal P_HR_NS71 : unsigned(11 downto 0);
	signal P_HR_NS72 : unsigned(11 downto 0);
	signal P_HR_NS73 : unsigned(11 downto 0);
	signal P_HR_NS74 : unsigned(11 downto 0);
	signal P_HR_NS75 : unsigned(11 downto 0);
	signal P_HR_NS76 : unsigned(11 downto 0);
	signal P_HR_NS77 : unsigned(11 downto 0);
	signal P_HR_NS78 : unsigned(11 downto 0);
	signal P_HR_NS79 : unsigned(11 downto 0);
	signal P_HR_NS80 : unsigned(11 downto 0);
	signal P_HR_NS81 : unsigned(11 downto 0);
	signal P_HR_NS82 : unsigned(11 downto 0);
	signal P_HR_NS83 : unsigned(11 downto 0);
	signal P_HR_NS84 : unsigned(11 downto 0);
	signal P_HR_NS85 : unsigned(11 downto 0);
	signal P_HR_NS86 : unsigned(11 downto 0);
	signal P_HR_NS87 : unsigned(11 downto 0);
	signal P_HR_NS88 : unsigned(11 downto 0);
	signal P_HR_NS89 : unsigned(11 downto 0);
	signal P_HR_NS90 : unsigned(11 downto 0);
	signal P_HR_NS91 : unsigned(11 downto 0);
	signal P_HR_NS92 : unsigned(11 downto 0);
	signal P_HR_NS93 : unsigned(11 downto 0);
	signal P_HR_NS94 : unsigned(11 downto 0);
	signal P_HR_NS95 : unsigned(11 downto 0);
	signal P_HR_NS96 : unsigned(11 downto 0);
	signal P_HR_NS97 : unsigned(11 downto 0);
	signal P_HR_NS98 : unsigned(11 downto 0);
	signal P_HR_NS99 : unsigned(11 downto 0);
	signal P_HR_NS100 : unsigned(11 downto 0);
	signal P_HR_NS101 : unsigned(11 downto 0);
	signal P_HR_NS102 : unsigned(11 downto 0);
	signal P_HR_NS103 : unsigned(11 downto 0);
	signal P_HR_NS104 : unsigned(11 downto 0);
	signal P_HR_NS105 : unsigned(11 downto 0);
	signal P_HR_NS106 : unsigned(11 downto 0);
	signal P_HR_NS107 : unsigned(11 downto 0);
	signal P_HR_NS108 : unsigned(11 downto 0);
	signal P_HR_NS109 : unsigned(11 downto 0);
	signal P_HR_NS110 : unsigned(11 downto 0);
	signal P_HR_NS111 : unsigned(11 downto 0);
	signal P_HR_NS112 : unsigned(11 downto 0);
	signal P_HR_NS113 : unsigned(11 downto 0);
	signal P_HR_NS114 : unsigned(11 downto 0);
	signal P_HR_NS115 : unsigned(11 downto 0);
	signal P_HR_NS116 : unsigned(11 downto 0);
	signal P_HR_NS117 : unsigned(11 downto 0);
	signal P_HR_NS118 : unsigned(11 downto 0);
	signal P_HR_NS119 : unsigned(11 downto 0);
	signal P_HR_NS120 : unsigned(11 downto 0);
	signal P_HR_NS121 : unsigned(11 downto 0);
	signal P_HR_NS122 : unsigned(11 downto 0);
	signal P_HR_NS123 : unsigned(11 downto 0);
	signal P_HR_NS124 : unsigned(11 downto 0);
	signal P_HR_NS125 : unsigned(11 downto 0);
	signal P_HR_NS126 : unsigned(11 downto 0);
	signal P_HR_NS127 : unsigned(11 downto 0);
	signal P_HR_NS128 : unsigned(11 downto 0);
	signal P_HR_NS129 : unsigned(11 downto 0);
	signal P_HR_NS130 : unsigned(11 downto 0);
	signal P_HR_NS131 : unsigned(11 downto 0);
	signal P_HR_NS132 : unsigned(11 downto 0);
	signal P_HR_NS133 : unsigned(11 downto 0);
	signal P_HR_NS134 : unsigned(11 downto 0);
	signal P_HR_NS135 : unsigned(11 downto 0);
	signal P_HR_NS136 : unsigned(11 downto 0);
	signal P_HR_NS137 : unsigned(11 downto 0);
	signal P_HR_NS138 : unsigned(11 downto 0);
	signal P_HR_NS139 : unsigned(11 downto 0);
	signal P_HR_NS140 : unsigned(11 downto 0);
	signal P_HR_NS141 : unsigned(11 downto 0);
	signal P_HR_NS142 : unsigned(11 downto 0);
	signal P_HR_NS143 : unsigned(11 downto 0);
	signal P_HR_NS144 : unsigned(11 downto 0);
	signal P_HR_NS145 : unsigned(11 downto 0);
	signal P_HR_NS146 : unsigned(11 downto 0);
	signal P_HR_NS147 : unsigned(11 downto 0);
	signal P_HR_NS148 : unsigned(11 downto 0);
	signal P_HR_NS149 : unsigned(11 downto 0);
	signal P_HR_NS150 : unsigned(11 downto 0);
	signal P_HR_NS151 : unsigned(11 downto 0);
	signal P_HR_NS152 : unsigned(11 downto 0);
	signal P_HR_NS153 : unsigned(11 downto 0);
	signal P_HR_NS154 : unsigned(11 downto 0);
	signal P_HR_NS155 : unsigned(11 downto 0);
	signal P_HR_NS156 : unsigned(11 downto 0);
	signal P_HR_NS157 : unsigned(11 downto 0);
	signal P_HR_NS158 : unsigned(11 downto 0);
	signal P_HR_NS159 : unsigned(11 downto 0);
	signal P_HR_NS160 : unsigned(11 downto 0);
	signal P_HR_NS161 : unsigned(11 downto 0);
	signal P_HR_NS162 : unsigned(11 downto 0);
	signal P_HR_NS163 : unsigned(11 downto 0);
	signal P_HR_NS164 : unsigned(11 downto 0);
	signal P_HR_NS165 : unsigned(11 downto 0);
	signal P_HR_NS166 : unsigned(11 downto 0);
	signal P_HR_NS167 : unsigned(11 downto 0);
	signal P_HR_NS168 : unsigned(11 downto 0);
	signal P_HR_NS169 : unsigned(11 downto 0);
	signal P_HR_NS170 : unsigned(11 downto 0);
	signal P_HR_NS171 : unsigned(11 downto 0);
	signal P_HR_NS172 : unsigned(11 downto 0);
	signal P_HR_NS173 : unsigned(11 downto 0);
	signal P_HR_NS174 : unsigned(11 downto 0);
	signal P_HR_NS175 : unsigned(11 downto 0);
	signal P_HR_NS176 : unsigned(11 downto 0);
	signal P_HR_NS177 : unsigned(11 downto 0);
	signal P_HR_NS178 : unsigned(11 downto 0);
	signal P_HR_NS179 : unsigned(11 downto 0);
	signal P_HR_NS180 : unsigned(11 downto 0);
	signal P_HR_NS181 : unsigned(11 downto 0);
	signal P_HR_NS182 : unsigned(11 downto 0);
	signal P_HR_NS183 : unsigned(11 downto 0);
	signal P_HR_NS184 : unsigned(11 downto 0);
	signal P_HR_NS185 : unsigned(11 downto 0);
	signal P_HR_NS186 : unsigned(11 downto 0);
	signal P_HR_NS187 : unsigned(11 downto 0);
	signal P_HR_NS188 : unsigned(11 downto 0);
	signal P_HR_NS189 : unsigned(11 downto 0);
	signal P_HR_NS190 : unsigned(11 downto 0);
	signal P_HR_NS191 : unsigned(11 downto 0);
	signal P_HR_NS192 : unsigned(11 downto 0);
	signal P_HR_NS193 : unsigned(11 downto 0);
	signal P_HR_NS194 : unsigned(11 downto 0);
	signal P_HR_NS195 : unsigned(11 downto 0);
	signal P_HR_NS196 : unsigned(11 downto 0);
	signal P_HR_NS197 : unsigned(11 downto 0);
	signal P_HR_NS198 : unsigned(11 downto 0);
	signal P_HR_NS199 : unsigned(11 downto 0);
	signal P_HR_NS200 : unsigned(11 downto 0);
	signal P_HR_NS201 : unsigned(11 downto 0);
	signal P_HR_NS202 : unsigned(11 downto 0);
	signal P_HR_NS203 : unsigned(11 downto 0);
	signal P_HR_NS204 : unsigned(11 downto 0);
	signal P_HR_NS205 : unsigned(11 downto 0);
	signal P_HR_NS206 : unsigned(11 downto 0);
	signal P_HR_NS207 : unsigned(11 downto 0);
	signal P_HR_NS208 : unsigned(11 downto 0);
	signal P_HR_NS209 : unsigned(11 downto 0);
	signal P_HR_NS210 : unsigned(11 downto 0);
	signal P_HR_NS211 : unsigned(11 downto 0);
	signal P_HR_NS212 : unsigned(11 downto 0);
	signal P_HR_NS213 : unsigned(11 downto 0);
	signal P_HR_NS214 : unsigned(11 downto 0);
	signal P_HR_NS215 : unsigned(11 downto 0);
	signal P_HR_NS216 : unsigned(11 downto 0);
	signal P_HR_NS217 : unsigned(11 downto 0);
	signal P_HR_NS218 : unsigned(11 downto 0);
	signal P_HR_NS219 : unsigned(11 downto 0);
	signal P_HR_NS220 : unsigned(11 downto 0);
	signal P_HR_NS221 : unsigned(11 downto 0);
	signal P_HR_NS222 : unsigned(11 downto 0);
	signal P_HR_NS223 : unsigned(11 downto 0);
	signal P_HR_NS224 : unsigned(11 downto 0);
	signal P_HR_NS225 : unsigned(11 downto 0);
	signal P_HR_NS226 : unsigned(11 downto 0);
	signal P_HR_NS227 : unsigned(11 downto 0);
	signal P_HR_NS228 : unsigned(11 downto 0);
	signal P_HR_NS229 : unsigned(11 downto 0);
	signal P_HR_NS230 : unsigned(11 downto 0);
	signal P_HR_NS231 : unsigned(11 downto 0);
	signal P_HR_NS232 : unsigned(11 downto 0);
	signal P_HR_NS233 : unsigned(11 downto 0);
	signal P_HR_NS234 : unsigned(11 downto 0);
	signal P_HR_NS235 : unsigned(11 downto 0);
	signal P_HR_NS236 : unsigned(11 downto 0);
	signal P_HR_NS237 : unsigned(11 downto 0);
	signal P_HR_NS238 : unsigned(11 downto 0);
	signal P_HR_NS239 : unsigned(11 downto 0);
	signal P_HR_NS240 : unsigned(11 downto 0);
	signal P_HR_NS241 : unsigned(11 downto 0);
	signal P_HR_NS242 : unsigned(11 downto 0);
	signal P_HR_NS243 : unsigned(11 downto 0);
	signal P_HR_NS244 : unsigned(11 downto 0);
	signal P_HR_NS245 : unsigned(11 downto 0);
	signal P_HR_NS246 : unsigned(11 downto 0);
	signal P_HR_NS247 : unsigned(11 downto 0);
	signal P_HR_NS248 : unsigned(11 downto 0);
	signal P_HR_NS249 : unsigned(11 downto 0);
	signal P_HR_NS250 : unsigned(11 downto 0);
	signal P_HR_NS251 : unsigned(11 downto 0);
	signal P_HR_NS252 : unsigned(11 downto 0);
	signal P_HR_NS253 : unsigned(11 downto 0);
	signal P_HR_NS254 : unsigned(11 downto 0);
	signal P_HR_NS255 : unsigned(11 downto 0);
	signal P_HR_NS256 : unsigned(11 downto 0);
	signal P_HR_NS257 : unsigned(11 downto 0);
	signal P_HR_NS258 : unsigned(11 downto 0);
	signal P_HR_NS259 : unsigned(11 downto 0);
	signal P_HR_NS260 : unsigned(11 downto 0);
	signal P_HR_NS261 : unsigned(11 downto 0);
	signal P_HR_NS262 : unsigned(11 downto 0);
	signal P_HR_NS263 : unsigned(11 downto 0);
	signal P_HR_NS264 : unsigned(11 downto 0);
	signal P_HR_NS265 : unsigned(11 downto 0);
	signal P_HR_NS266 : unsigned(11 downto 0);
	signal P_HR_NS267 : unsigned(11 downto 0);
	signal P_HR_NS268 : unsigned(11 downto 0);
	signal P_HR_NS269 : unsigned(11 downto 0);
	signal P_HR_NS270 : unsigned(11 downto 0);
	signal P_HR_NS271 : unsigned(11 downto 0);
	signal P_HR_NS272 : unsigned(11 downto 0);
	signal P_HR_NS273 : unsigned(11 downto 0);
	signal P_HR_NS274 : unsigned(11 downto 0);
	signal P_HR_NS275 : unsigned(11 downto 0);
	signal P_HR_NS276 : unsigned(11 downto 0);
	signal P_HR_NS277 : unsigned(11 downto 0);
	signal P_HR_NS278 : unsigned(11 downto 0);
	signal P_HR_NS279 : unsigned(11 downto 0);
	signal P_HR_NS280 : unsigned(11 downto 0);
	signal P_HR_NS281 : unsigned(11 downto 0);
	signal P_HR_NS282 : unsigned(11 downto 0);
	signal P_HR_NS283 : unsigned(11 downto 0);
	signal P_HR_NS284 : unsigned(11 downto 0);
	signal P_HR_NS285 : unsigned(11 downto 0);
	signal P_HR_NS286 : unsigned(11 downto 0);
	signal P_HR_NS287 : unsigned(11 downto 0);
	signal P_HR_NS288 : unsigned(11 downto 0);
	signal P_HR_NS289 : unsigned(11 downto 0);
	signal P_HR_NS290 : unsigned(11 downto 0);
	signal P_HR_NS291 : unsigned(11 downto 0);
	signal P_HR_NS292 : unsigned(11 downto 0);
	signal P_HR_NS293 : unsigned(11 downto 0);
	signal P_HR_NS294 : unsigned(11 downto 0);
	signal P_HR_NS295 : unsigned(11 downto 0);
	signal P_HR_NS296 : unsigned(11 downto 0);
	signal P_HR_NS297 : unsigned(11 downto 0);
	signal P_HR_NS298 : unsigned(11 downto 0);
	signal P_HR_NS299 : unsigned(11 downto 0);
	signal P_HR_NS300 : unsigned(11 downto 0);
	signal P_HR_NS301 : unsigned(11 downto 0);
	signal P_HR_NS302 : unsigned(11 downto 0);
	signal P_HR_NS303 : unsigned(11 downto 0);
	signal P_HR_NS304 : unsigned(11 downto 0);
	signal P_HR_NS305 : unsigned(11 downto 0);
	signal P_HR_NS306 : unsigned(11 downto 0);
	signal P_HR_NS307 : unsigned(11 downto 0);
	signal P_HR_NS308 : unsigned(11 downto 0);
	signal P_HR_NS309 : unsigned(11 downto 0);
	signal P_HR_NS310 : unsigned(11 downto 0);
	signal P_HR_NS311 : unsigned(11 downto 0);
	signal P_HR_NS312 : unsigned(11 downto 0);
	signal P_HR_NS313 : unsigned(11 downto 0);
	signal P_HR_NS314 : unsigned(11 downto 0);
	signal P_HR_NS315 : unsigned(11 downto 0);
	signal P_HR_NS316 : unsigned(11 downto 0);
	signal P_HR_NS317 : unsigned(11 downto 0);
	signal P_HR_NS318 : unsigned(11 downto 0);
	signal P_HR_NS319 : unsigned(11 downto 0);
	signal P_HR_NS320 : unsigned(11 downto 0);
	signal P_HR_NS321 : unsigned(11 downto 0);
	signal P_HR_NS322 : unsigned(11 downto 0);
	signal P_HR_NS323 : unsigned(11 downto 0);
	signal P_HR_NS324 : unsigned(11 downto 0);
	signal P_HR_NS325 : unsigned(11 downto 0);
	signal P_HR_NS326 : unsigned(11 downto 0);
	signal P_HR_NS327 : unsigned(11 downto 0);
	signal P_HR_NS328 : unsigned(11 downto 0);
	signal P_HR_NS329 : unsigned(11 downto 0);
	signal P_HR_NS330 : unsigned(11 downto 0);
	signal P_HR_NS331 : unsigned(11 downto 0);
	signal P_HR_NS332 : unsigned(11 downto 0);
	signal P_HR_NS333 : unsigned(11 downto 0);
	signal P_HR_NS334 : unsigned(11 downto 0);
	signal P_HR_NS335 : unsigned(11 downto 0);
	signal P_HR_NS336 : unsigned(11 downto 0);
	signal P_HR_NS337 : unsigned(11 downto 0);
	signal P_HR_NS338 : unsigned(11 downto 0);
	signal P_HR_NS339 : unsigned(11 downto 0);
	signal P_HR_NS340 : unsigned(11 downto 0);
	signal P_HR_NS341 : unsigned(11 downto 0);
	signal P_HR_NS342 : unsigned(11 downto 0);
	signal P_HR_NS343 : unsigned(11 downto 0);
	signal P_HR_NS344 : unsigned(11 downto 0);
	signal P_HR_NS345 : unsigned(11 downto 0);
	signal P_HR_NS346 : unsigned(11 downto 0);
	signal P_HR_NS347 : unsigned(11 downto 0);
	signal P_HR_NS348 : unsigned(11 downto 0);
	signal P_HR_NS349 : unsigned(11 downto 0);
	signal P_HR_NS350 : unsigned(11 downto 0);
	signal P_HR_NS351 : unsigned(11 downto 0);
	signal P_HR_NS352 : unsigned(11 downto 0);
	signal P_HR_NS353 : unsigned(11 downto 0);
	signal P_HR_NS354 : unsigned(11 downto 0);
	signal P_HR_NS355 : unsigned(11 downto 0);
	signal P_HR_NS356 : unsigned(11 downto 0);
	signal P_HR_NS357 : unsigned(11 downto 0);
	signal P_HR_NS358 : unsigned(11 downto 0);
	signal P_HR_NS359 : unsigned(11 downto 0);
	signal P_HR_NS360 : unsigned(11 downto 0);
	signal P_HR_NS361 : unsigned(11 downto 0);
	signal P_HR_NS362 : unsigned(11 downto 0);
	signal P_HR_NS363 : unsigned(11 downto 0);
	signal P_HR_NS364 : unsigned(11 downto 0);
	signal P_HR_NS365 : unsigned(11 downto 0);
	signal P_HR_NS366 : unsigned(11 downto 0);
	signal P_HR_NS367 : unsigned(11 downto 0);
	signal P_HR_NS368 : unsigned(11 downto 0);
	signal P_HR_NS369 : unsigned(11 downto 0);
	signal P_HR_NS370 : unsigned(11 downto 0);
	signal P_HR_NS371 : unsigned(11 downto 0);
	signal P_HR_NS372 : unsigned(11 downto 0);
	signal P_HR_NS373 : unsigned(11 downto 0);
	signal P_HR_NS374 : unsigned(11 downto 0);
	signal P_HR_NS375 : unsigned(11 downto 0);
	signal P_HR_NS376 : unsigned(11 downto 0);
	signal P_HR_NS377 : unsigned(11 downto 0);
	signal P_HR_NS378 : unsigned(11 downto 0);
	signal P_HR_NS379 : unsigned(11 downto 0);
	signal P_HR_NS380 : unsigned(11 downto 0);
	signal P_HR_NS381 : unsigned(11 downto 0);
	signal P_HR_NS382 : unsigned(11 downto 0);
	signal P_HR_NS383 : unsigned(11 downto 0);
	signal P_HR_NS384 : unsigned(11 downto 0);
	signal P_HR_NS385 : unsigned(11 downto 0);
	signal P_HR_NS386 : unsigned(11 downto 0);
	signal P_HR_NS387 : unsigned(11 downto 0);
	signal P_HR_NS388 : unsigned(11 downto 0);
	signal P_HR_NS389 : unsigned(11 downto 0);
	signal P_HR_NS390 : unsigned(11 downto 0);
	signal P_HR_NS391 : unsigned(11 downto 0);
	signal P_HR_NS392 : unsigned(11 downto 0);
	signal P_HR_NS393 : unsigned(11 downto 0);
	signal P_HR_NS394 : unsigned(11 downto 0);
	signal P_HR_NS395 : unsigned(11 downto 0);
	signal P_HR_NS396 : unsigned(11 downto 0);
	signal P_HR_NS397 : unsigned(11 downto 0);
	signal P_HR_NS398 : unsigned(11 downto 0);
	signal P_HR_NS399 : unsigned(11 downto 0);
	signal P_HR_NS400 : unsigned(11 downto 0);
	signal P_HR_NS401 : unsigned(11 downto 0);
	signal P_HR_NS402 : unsigned(11 downto 0);
	signal P_HR_NS403 : unsigned(11 downto 0);
	signal P_HR_NS404 : unsigned(11 downto 0);
	signal P_HR_NS405 : unsigned(11 downto 0);
	signal P_HR_NS406 : unsigned(11 downto 0);
	signal P_HR_NS407 : unsigned(11 downto 0);
	signal P_HR_NS408 : unsigned(11 downto 0);
	signal P_HR_NS409 : unsigned(11 downto 0);
	signal P_HR_NS410 : unsigned(11 downto 0);
	signal P_HR_NS411 : unsigned(11 downto 0);
	signal P_HR_NS412 : unsigned(11 downto 0);
	signal P_HR_NS413 : unsigned(11 downto 0);
	signal P_HR_NS414 : unsigned(11 downto 0);
	signal P_HR_NS415 : unsigned(11 downto 0);
	signal P_HR_NS416 : unsigned(11 downto 0);
	signal P_HR_NS417 : unsigned(11 downto 0);
	signal P_HR_NS418 : unsigned(11 downto 0);
	signal P_HR_NS419 : unsigned(11 downto 0);
	signal P_HR_NS420 : unsigned(11 downto 0);
	signal P_HR_NS421 : unsigned(11 downto 0);
	signal P_HR_NS422 : unsigned(11 downto 0);
	signal P_HR_NS423 : unsigned(11 downto 0);
	signal P_HR_NS424 : unsigned(11 downto 0);
	signal P_HR_NS425 : unsigned(11 downto 0);
	signal P_HR_NS426 : unsigned(11 downto 0);
	signal P_HR_NS427 : unsigned(11 downto 0);
	signal P_HR_NS428 : unsigned(11 downto 0);
	signal P_HR_NS429 : unsigned(11 downto 0);
	signal P_HR_NS430 : unsigned(11 downto 0);
	signal P_HR_NS431 : unsigned(11 downto 0);
	signal P_HR_NS432 : unsigned(11 downto 0);
	signal P_HR_NS433 : unsigned(11 downto 0);
	signal P_HR_NS434 : unsigned(11 downto 0);
	signal P_HR_NS435 : unsigned(11 downto 0);
	signal P_HR_NS436 : unsigned(11 downto 0);
	signal P_HR_NS437 : unsigned(11 downto 0);
	signal P_HR_NS438 : unsigned(11 downto 0);
	signal P_HR_NS439 : unsigned(11 downto 0);
	signal P_HR_NS440 : unsigned(11 downto 0);
	signal P_HR_NS441 : unsigned(11 downto 0);
	signal P_HR_NS442 : unsigned(11 downto 0);
	signal P_HR_NS443 : unsigned(11 downto 0);
	signal P_HR_NS444 : unsigned(11 downto 0);
	signal P_HR_NS445 : unsigned(11 downto 0);
	signal P_HR_NS446 : unsigned(11 downto 0);
	signal P_HR_NS447 : unsigned(11 downto 0);
	signal P_HR_NS448 : unsigned(11 downto 0);
	signal P_HR_NS449 : unsigned(11 downto 0);
	signal P_HR_NS450 : unsigned(11 downto 0);
	signal P_HR_NS451 : unsigned(11 downto 0);
	signal P_HR_NS452 : unsigned(11 downto 0);
	signal P_HR_NS453 : unsigned(11 downto 0);
	signal P_HR_NS454 : unsigned(11 downto 0);
	signal P_HR_NS455 : unsigned(11 downto 0);
	signal P_HR_NS456 : unsigned(11 downto 0);
	signal P_HR_NS457 : unsigned(11 downto 0);
	signal P_HR_NS458 : unsigned(11 downto 0);
		
	signal P_EDA_NS1 : unsigned(11 downto 0);
	signal P_EDA_NS2 : unsigned(11 downto 0);
	signal P_EDA_NS3 : unsigned(11 downto 0);
	signal P_EDA_NS4 : unsigned(11 downto 0);
	signal P_EDA_NS5 : unsigned(11 downto 0);
	signal P_EDA_NS6 : unsigned(11 downto 0);
	signal P_EDA_NS7 : unsigned(11 downto 0);
	signal P_EDA_NS8 : unsigned(11 downto 0);
	signal P_EDA_NS9 : unsigned(11 downto 0);
	signal P_EDA_NS10 : unsigned(11 downto 0);
	signal P_EDA_NS11 : unsigned(11 downto 0);
	signal P_EDA_NS12 : unsigned(11 downto 0);
	signal P_EDA_NS13 : unsigned(11 downto 0);
	signal P_EDA_NS14 : unsigned(11 downto 0);
	signal P_EDA_NS15 : unsigned(11 downto 0);
	signal P_EDA_NS16 : unsigned(11 downto 0);
	signal P_EDA_NS17 : unsigned(11 downto 0);
	signal P_EDA_NS18 : unsigned(11 downto 0);
	signal P_EDA_NS19 : unsigned(11 downto 0);
	signal P_EDA_NS20 : unsigned(11 downto 0);
	signal P_EDA_NS21 : unsigned(11 downto 0);
	signal P_EDA_NS22 : unsigned(11 downto 0);
	signal P_EDA_NS23 : unsigned(11 downto 0);
	signal P_EDA_NS24 : unsigned(11 downto 0);
	signal P_EDA_NS25 : unsigned(11 downto 0);
	signal P_EDA_NS26 : unsigned(11 downto 0);
	signal P_EDA_NS27 : unsigned(11 downto 0);
	signal P_EDA_NS28 : unsigned(11 downto 0);
	signal P_EDA_NS29 : unsigned(11 downto 0);
	signal P_EDA_NS30 : unsigned(11 downto 0);
	signal P_EDA_NS31 : unsigned(11 downto 0);
	signal P_EDA_NS32 : unsigned(11 downto 0);
	signal P_EDA_NS33 : unsigned(11 downto 0);
	signal P_EDA_NS34 : unsigned(11 downto 0);
	signal P_EDA_NS35 : unsigned(11 downto 0);
	signal P_EDA_NS36 : unsigned(11 downto 0);
	signal P_EDA_NS37 : unsigned(11 downto 0);
	signal P_EDA_NS38 : unsigned(11 downto 0);
	signal P_EDA_NS39 : unsigned(11 downto 0);
	signal P_EDA_NS40 : unsigned(11 downto 0);
	signal P_EDA_NS41 : unsigned(11 downto 0);
	signal P_EDA_NS42 : unsigned(11 downto 0);
	signal P_EDA_NS43 : unsigned(11 downto 0);
	signal P_EDA_NS44 : unsigned(11 downto 0);
	signal P_EDA_NS45 : unsigned(11 downto 0);
	signal P_EDA_NS46 : unsigned(11 downto 0);
	signal P_EDA_NS47 : unsigned(11 downto 0);
	signal P_EDA_NS48 : unsigned(11 downto 0);
	signal P_EDA_NS49 : unsigned(11 downto 0);
	signal P_EDA_NS50 : unsigned(11 downto 0);
	signal P_EDA_NS51 : unsigned(11 downto 0);
	signal P_EDA_NS52 : unsigned(11 downto 0);
	signal P_EDA_NS53 : unsigned(11 downto 0);
	signal P_EDA_NS54 : unsigned(11 downto 0);
	signal P_EDA_NS55 : unsigned(11 downto 0);
	signal P_EDA_NS56 : unsigned(11 downto 0);
	signal P_EDA_NS57 : unsigned(11 downto 0);
	signal P_EDA_NS58 : unsigned(11 downto 0);
	signal P_EDA_NS59 : unsigned(11 downto 0);
	signal P_EDA_NS60 : unsigned(11 downto 0);
	signal P_EDA_NS61 : unsigned(11 downto 0);
	signal P_EDA_NS62 : unsigned(11 downto 0);
	signal P_EDA_NS63 : unsigned(11 downto 0);
	signal P_EDA_NS64 : unsigned(11 downto 0);
	signal P_EDA_NS65 : unsigned(11 downto 0);
	signal P_EDA_NS66 : unsigned(11 downto 0);
	signal P_EDA_NS67 : unsigned(11 downto 0);
	
	signal P_TEMP_S : unsigned(11 downto 0);
	signal P_TEMP_NS : unsigned(11 downto 0);
	
	signal P_EDA_S : unsigned(11 downto 0);
	signal P_EDA_NS : unsigned(11 downto 0);
	
	signal P_HR_S : unsigned(11 downto 0);
	signal P_HR_NS : unsigned(11 downto 0);
	
	signal stress_score : unsigned(47 downto 0);
	signal not_stress_score : unsigned(48 downto 0);
	
	type type_state is (NORMAL, TRAINING_S, TRAINING_NS);
	attribute enum_encoding : string;
	attribute enum_encoding of type_state : type is "00 01 11";
	
	signal state, next_state: type_state;
	
	-- constants
    constant P_STRESS : unsigned(11 downto 0) := "011111010000"; -- 20
	constant P_NOT_STRESS : unsigned(12 downto 0) := "1111101000000"; -- 80
	
	--constant P_STRESS : unsigned(12 downto 0) := "1001110001000"; 
	--constant P_NOT_STRESS : unsigned(12 downto 0) := "1001110001000";
	
begin
	
	process(clk, rst) --state transition
	begin
		if (rst = '1') then
			state <= NORMAL;
		elsif (rising_edge(clk)) then
			state <= next_state;
		end if;
	end process;
	
	process(state, s1) -- combinational state assignment
	begin
		case state is
			when NORMAL =>
				if s1 = "01" then
					next_state <= TRAINING_S;
				elsif s1 = "11" then
					next_state <= TRAINING_NS;
				else
					next_state <= NORMAL;
				end if;
			when TRAINING_S =>
				if s1 = "01" then
					next_state <= TRAINING_S;
				elsif s1 = "11" then
					next_state <= TRAINING_NS;
				else
					next_state <= NORMAL;
				end if;
			when TRAINING_NS =>
				if s1 = "01" then
					next_state <= TRAINING_S;
				elsif s1 = "11" then
					next_state <= TRAINING_NS;
				else
					next_state <= NORMAL;
				end if;
			when others => null;
		end case;
	end process;
	
	-- should expect status = 11 when in training mode
	process(clk,rst) -- output block
	begin
		if (rst = '1') then
			status <= "00";
		elsif (rising_edge(clk)) then
			if stress_score < not_stress_score then
				status <= "01"; -- not stressed
			elsif stress_score > not_stress_score then
				status <= "10"; -- stressed
			elsif stress_score = not_stress_score then
				status <= "11"; -- rare, equality
			else
				status <= "00";
			end if;

		end if;	
	end process;	
	

	process(clk, rst) -- stress score
	begin
		if (rst = '1') then
		-- reset logic
		P_TEMP_S1 <= (others => '0');
		P_TEMP_S2 <= (others => '0');
		P_TEMP_S3 <= (others => '0');
		P_TEMP_S4 <= (others => '0');
		P_TEMP_S5 <= (others => '0');
		P_TEMP_S6 <= (others => '0');
		P_TEMP_S7 <= (others => '0');
		P_TEMP_S8 <= (others => '0');
		P_TEMP_S9 <= (others => '0');
		P_TEMP_S10 <= (others => '0');
		P_TEMP_S11 <= (others => '0');
		P_TEMP_S12 <= (others => '0');
		P_TEMP_S13 <= (others => '0');
		P_TEMP_S14 <= (others => '0');
		P_TEMP_S15 <= (others => '0');
		P_TEMP_S16 <= (others => '0');
		P_TEMP_S17 <= (others => '0');
		P_TEMP_S18 <= (others => '0');
		P_TEMP_S19 <= (others => '0');
		P_TEMP_S20 <= (others => '0');
		P_TEMP_S21 <= (others => '0');
		P_TEMP_S22 <= (others => '0');
		P_TEMP_S23 <= (others => '0');
		P_TEMP_S24 <= (others => '0');
		P_TEMP_S25 <= (others => '0');
		P_TEMP_S26 <= (others => '0');
		P_TEMP_S27 <= (others => '0');
		P_TEMP_S28 <= (others => '0');
		P_TEMP_S29 <= (others => '0');
		P_TEMP_S30 <= (others => '0');
			
		P_EDA_S1 <= (others => '0');
		P_EDA_S2 <= (others => '0');
		P_EDA_S3 <= (others => '0');
		P_EDA_S4 <= (others => '0');
		P_EDA_S5 <= (others => '0');
		P_EDA_S6 <= (others => '0');
		P_EDA_S7 <= (others => '0');
		P_EDA_S8 <= (others => '0');
		P_EDA_S9 <= (others => '0');
		P_EDA_S10 <= (others => '0');
		P_EDA_S11 <= (others => '0');
		P_EDA_S12 <= (others => '0');
		P_EDA_S13 <= (others => '0');
		P_EDA_S14 <= (others => '0');
		P_EDA_S15 <= (others => '0');
		P_EDA_S16 <= (others => '0');
		P_EDA_S17 <= (others => '0');
		P_EDA_S18 <= (others => '0');
		P_EDA_S19 <= (others => '0');
		P_EDA_S20 <= (others => '0');
		P_EDA_S21 <= (others => '0');
		P_EDA_S22 <= (others => '0');
		P_EDA_S23 <= (others => '0');
		P_EDA_S24 <= (others => '0');
		P_EDA_S25 <= (others => '0');
		P_EDA_S26 <= (others => '0');
		P_EDA_S27 <= (others => '0');
		P_EDA_S28 <= (others => '0');
		P_EDA_S29 <= (others => '0');
		P_EDA_S30 <= (others => '0');
		P_EDA_S31 <= (others => '0');
		P_EDA_S32 <= (others => '0');
		P_EDA_S33 <= (others => '0');
		P_EDA_S34 <= (others => '0');
		P_EDA_S35 <= (others => '0');
		P_EDA_S36 <= (others => '0');
		P_EDA_S37 <= (others => '0');
		P_EDA_S38 <= (others => '0');
		P_EDA_S39 <= (others => '0');
		P_EDA_S40 <= (others => '0');
		P_EDA_S41 <= (others => '0');
		P_EDA_S42 <= (others => '0');
		P_EDA_S43 <= (others => '0');
		P_EDA_S44 <= (others => '0');
		P_EDA_S45 <= (others => '0');
		P_EDA_S46 <= (others => '0');
		P_EDA_S47 <= (others => '0');
		P_EDA_S48 <= (others => '0');
		P_EDA_S49 <= (others => '0');
		P_EDA_S50 <= (others => '0');
		P_EDA_S51 <= (others => '0');
		P_EDA_S52 <= (others => '0');
		P_EDA_S53 <= (others => '0');
		P_EDA_S54 <= (others => '0');
		P_EDA_S55 <= (others => '0');
		P_EDA_S56 <= (others => '0');
		P_EDA_S57 <= (others => '0');
		P_EDA_S58 <= (others => '0');
		P_EDA_S59 <= (others => '0');
		P_EDA_S60 <= (others => '0');
		P_EDA_S61 <= (others => '0');
		P_EDA_S62 <= (others => '0');
		P_EDA_S63 <= (others => '0');
		P_EDA_S64 <= (others => '0');
		P_EDA_S65 <= (others => '0');	
			
		P_HR_S1 <= (others => '0');
		P_HR_S2 <= (others => '0');
		P_HR_S3 <= (others => '0');
		P_HR_S4 <= (others => '0');
		P_HR_S5 <= (others => '0');
		P_HR_S6 <= (others => '0');
		P_HR_S7 <= (others => '0');
		P_HR_S8 <= (others => '0');
		P_HR_S9 <= (others => '0');
		P_HR_S10 <= (others => '0');
		P_HR_S11 <= (others => '0');
		P_HR_S12 <= (others => '0');
		P_HR_S13 <= (others => '0');
		P_HR_S14 <= (others => '0');
		P_HR_S15 <= (others => '0');
		P_HR_S16 <= (others => '0');
		P_HR_S17 <= (others => '0');
		P_HR_S18 <= (others => '0');
		P_HR_S19 <= (others => '0');
		P_HR_S20 <= (others => '0');
		P_HR_S21 <= (others => '0');
		P_HR_S22 <= (others => '0');
		P_HR_S23 <= (others => '0');
		P_HR_S24 <= (others => '0');
		P_HR_S25 <= (others => '0');
		P_HR_S26 <= (others => '0');
		P_HR_S27 <= (others => '0');
		P_HR_S28 <= (others => '0');
		P_HR_S29 <= (others => '0');
		P_HR_S30 <= (others => '0');
		P_HR_S31 <= (others => '0');
		P_HR_S32 <= (others => '0');
		P_HR_S33 <= (others => '0');
		P_HR_S34 <= (others => '0');
		P_HR_S35 <= (others => '0');
		P_HR_S36 <= (others => '0');
		P_HR_S37 <= (others => '0');
		P_HR_S38 <= (others => '0');
		P_HR_S39 <= (others => '0');
		P_HR_S40 <= (others => '0');
		P_HR_S41 <= (others => '0');
		P_HR_S42 <= (others => '0');
		P_HR_S43 <= (others => '0');
		P_HR_S44 <= (others => '0');
		P_HR_S45 <= (others => '0');
		P_HR_S46 <= (others => '0');
		P_HR_S47 <= (others => '0');
		P_HR_S48 <= (others => '0');
		P_HR_S49 <= (others => '0');
		P_HR_S50 <= (others => '0');
		P_HR_S51 <= (others => '0');
		P_HR_S52 <= (others => '0');
		P_HR_S53 <= (others => '0');
		P_HR_S54 <= (others => '0');
		P_HR_S55 <= (others => '0');
		P_HR_S56 <= (others => '0');
		P_HR_S57 <= (others => '0');
		P_HR_S58 <= (others => '0');
		P_HR_S59 <= (others => '0');
		P_HR_S60 <= (others => '0');
		P_HR_S61 <= (others => '0');
		P_HR_S62 <= (others => '0');
		P_HR_S63 <= (others => '0');
		P_HR_S64 <= (others => '0');
		P_HR_S65 <= (others => '0');
		P_HR_S66 <= (others => '0');
		P_HR_S67 <= (others => '0');
		P_HR_S68 <= (others => '0');
		P_HR_S69 <= (others => '0');
		P_HR_S70 <= (others => '0');
		P_HR_S71 <= (others => '0');
		P_HR_S72 <= (others => '0');
		P_HR_S73 <= (others => '0');
		P_HR_S74 <= (others => '0');
		P_HR_S75 <= (others => '0');
		P_HR_S76 <= (others => '0');
		P_HR_S77 <= (others => '0');
		P_HR_S78 <= (others => '0');
		P_HR_S79 <= (others => '0');
		P_HR_S80 <= (others => '0');
		P_HR_S81 <= (others => '0');
		P_HR_S82 <= (others => '0');
		P_HR_S83 <= (others => '0');
		P_HR_S84 <= (others => '0');
		P_HR_S85 <= (others => '0');
		P_HR_S86 <= (others => '0');
		P_HR_S87 <= (others => '0');
		P_HR_S88 <= (others => '0');
		P_HR_S89 <= (others => '0');
		P_HR_S90 <= (others => '0');
		P_HR_S91 <= (others => '0');
		P_HR_S92 <= (others => '0');
		P_HR_S93 <= (others => '0');
		P_HR_S94 <= (others => '0');
		P_HR_S95 <= (others => '0');
		P_HR_S96 <= (others => '0');
		P_HR_S97 <= (others => '0');
		P_HR_S98 <= (others => '0');
		P_HR_S99 <= (others => '0');
		P_HR_S100 <= (others => '0');
		P_HR_S101 <= (others => '0');
		P_HR_S102 <= (others => '0');
		P_HR_S103 <= (others => '0');
		P_HR_S104 <= (others => '0');
		P_HR_S105 <= (others => '0');
		P_HR_S106 <= (others => '0');
		P_HR_S107 <= (others => '0');
		P_HR_S108 <= (others => '0');
		P_HR_S109 <= (others => '0');
		P_HR_S110 <= (others => '0');
		P_HR_S111 <= (others => '0');
		P_HR_S112 <= (others => '0');
		P_HR_S113 <= (others => '0');
		P_HR_S114 <= (others => '0');
		P_HR_S115 <= (others => '0');
		P_HR_S116 <= (others => '0');
		P_HR_S117 <= (others => '0');
		P_HR_S118 <= (others => '0');
		P_HR_S119 <= (others => '0');
		P_HR_S120 <= (others => '0');
		P_HR_S121 <= (others => '0');
		P_HR_S122 <= (others => '0');
		P_HR_S123 <= (others => '0');
		P_HR_S124 <= (others => '0');
		P_HR_S125 <= (others => '0');
		P_HR_S126 <= (others => '0');
		P_HR_S127 <= (others => '0');
		P_HR_S128 <= (others => '0');
		P_HR_S129 <= (others => '0');
		P_HR_S130 <= (others => '0');
		P_HR_S131 <= (others => '0');
		P_HR_S132 <= (others => '0');
		P_HR_S133 <= (others => '0');
		P_HR_S134 <= (others => '0');
		P_HR_S135 <= (others => '0');
		P_HR_S136 <= (others => '0');
		P_HR_S137 <= (others => '0');
		P_HR_S138 <= (others => '0');
		P_HR_S139 <= (others => '0');
		P_HR_S140 <= (others => '0');
		P_HR_S141 <= (others => '0');
		P_HR_S142 <= (others => '0');
		P_HR_S143 <= (others => '0');
		P_HR_S144 <= (others => '0');
		P_HR_S145 <= (others => '0');
		P_HR_S146 <= (others => '0');
		P_HR_S147 <= (others => '0');
		P_HR_S148 <= (others => '0');
		P_HR_S149 <= (others => '0');
		P_HR_S150 <= (others => '0');
		P_HR_S151 <= (others => '0');
		P_HR_S152 <= (others => '0');
		P_HR_S153 <= (others => '0');
		P_HR_S154 <= (others => '0');
		P_HR_S155 <= (others => '0');
		P_HR_S156 <= (others => '0');
		P_HR_S157 <= (others => '0');
		P_HR_S158 <= (others => '0');
		P_HR_S159 <= (others => '0');
		P_HR_S160 <= (others => '0');
		P_HR_S161 <= (others => '0');
		P_HR_S162 <= (others => '0');
		P_HR_S163 <= (others => '0');
		P_HR_S164 <= (others => '0');
		P_HR_S165 <= (others => '0');
		P_HR_S166 <= (others => '0');
		P_HR_S167 <= (others => '0');
		P_HR_S168 <= (others => '0');
		P_HR_S169 <= (others => '0');
		P_HR_S170 <= (others => '0');
		P_HR_S171 <= (others => '0');
		P_HR_S172 <= (others => '0');
		P_HR_S173 <= (others => '0');
		P_HR_S174 <= (others => '0');
		P_HR_S175 <= (others => '0');
		P_HR_S176 <= (others => '0');
		P_HR_S177 <= (others => '0');
		P_HR_S178 <= (others => '0');
		P_HR_S179 <= (others => '0');
		P_HR_S180 <= (others => '0');
		P_HR_S181 <= (others => '0');
		P_HR_S182 <= (others => '0');
		P_HR_S183 <= (others => '0');
		P_HR_S184 <= (others => '0');
		P_HR_S185 <= (others => '0');
		P_HR_S186 <= (others => '0');
		P_HR_S187 <= (others => '0');
		P_HR_S188 <= (others => '0');
		P_HR_S189 <= (others => '0');
		P_HR_S190 <= (others => '0');
		P_HR_S191 <= (others => '0');
		P_HR_S192 <= (others => '0');
		P_HR_S193 <= (others => '0');
		P_HR_S194 <= (others => '0');
		P_HR_S195 <= (others => '0');
		P_HR_S196 <= (others => '0');
		P_HR_S197 <= (others => '0');
		P_HR_S198 <= (others => '0');
		P_HR_S199 <= (others => '0');
		P_HR_S200 <= (others => '0');
		P_HR_S201 <= (others => '0');
		P_HR_S202 <= (others => '0');
		P_HR_S203 <= (others => '0');
		P_HR_S204 <= (others => '0');
		P_HR_S205 <= (others => '0');
		P_HR_S206 <= (others => '0');
		P_HR_S207 <= (others => '0');
		P_HR_S208 <= (others => '0');
		P_HR_S209 <= (others => '0');
		P_HR_S210 <= (others => '0');
		P_HR_S211 <= (others => '0');
		P_HR_S212 <= (others => '0');
		P_HR_S213 <= (others => '0');
		P_HR_S214 <= (others => '0');
		P_HR_S215 <= (others => '0');
		P_HR_S216 <= (others => '0');
		P_HR_S217 <= (others => '0');
		P_HR_S218 <= (others => '0');
		P_HR_S219 <= (others => '0');
		P_HR_S220 <= (others => '0');
		P_HR_S221 <= (others => '0');
		P_HR_S222 <= (others => '0');
		P_HR_S223 <= (others => '0');
		P_HR_S224 <= (others => '0');
		P_HR_S225 <= (others => '0');
		P_HR_S226 <= (others => '0');
		P_HR_S227 <= (others => '0');
		P_HR_S228 <= (others => '0');
		P_HR_S229 <= (others => '0');
		P_HR_S230 <= (others => '0');
		P_HR_S231 <= (others => '0');
		P_HR_S232 <= (others => '0');
		P_HR_S233 <= (others => '0');
		P_HR_S234 <= (others => '0');
		P_HR_S235 <= (others => '0');
		P_HR_S236 <= (others => '0');
		P_HR_S237 <= (others => '0');
		P_HR_S238 <= (others => '0');
		P_HR_S239 <= (others => '0');
		P_HR_S240 <= (others => '0');
		P_HR_S241 <= (others => '0');
		P_HR_S242 <= (others => '0');
		P_HR_S243 <= (others => '0');
		P_HR_S244 <= (others => '0');
		P_HR_S245 <= (others => '0');
		P_HR_S246 <= (others => '0');
		P_HR_S247 <= (others => '0');
		P_HR_S248 <= (others => '0');
		P_HR_S249 <= (others => '0');
		P_HR_S250 <= (others => '0');
		P_HR_S251 <= (others => '0');
		P_HR_S252 <= (others => '0');
		P_HR_S253 <= (others => '0');
		P_HR_S254 <= (others => '0');
		P_HR_S255 <= (others => '0');
		P_HR_S256 <= (others => '0');
		P_HR_S257 <= (others => '0');
		P_HR_S258 <= (others => '0');
		P_HR_S259 <= (others => '0');
		P_HR_S260 <= (others => '0');
		P_HR_S261 <= (others => '0');
		P_HR_S262 <= (others => '0');
		P_HR_S263 <= (others => '0');
		P_HR_S264 <= (others => '0');
		P_HR_S265 <= (others => '0');
		P_HR_S266 <= (others => '0');
		P_HR_S267 <= (others => '0');
		P_HR_S268 <= (others => '0');
		P_HR_S269 <= (others => '0');
		P_HR_S270 <= (others => '0');
		P_HR_S271 <= (others => '0');
		P_HR_S272 <= (others => '0');
		P_HR_S273 <= (others => '0');
		P_HR_S274 <= (others => '0');
		P_HR_S275 <= (others => '0');
		P_HR_S276 <= (others => '0');
		P_HR_S277 <= (others => '0');
		P_HR_S278 <= (others => '0');
		P_HR_S279 <= (others => '0');
		P_HR_S280 <= (others => '0');
		P_HR_S281 <= (others => '0');
		P_HR_S282 <= (others => '0');
		P_HR_S283 <= (others => '0');
		P_HR_S284 <= (others => '0');
		P_HR_S285 <= (others => '0');
		P_HR_S286 <= (others => '0');
		P_HR_S287 <= (others => '0');
		P_HR_S288 <= (others => '0');
		P_HR_S289 <= (others => '0');
		P_HR_S290 <= (others => '0');
		P_HR_S291 <= (others => '0');
		P_HR_S292 <= (others => '0');
		P_HR_S293 <= (others => '0');
		P_HR_S294 <= (others => '0');
		P_HR_S295 <= (others => '0');
		P_HR_S296 <= (others => '0');
		P_HR_S297 <= (others => '0');
		P_HR_S298 <= (others => '0');
		P_HR_S299 <= (others => '0');
		P_HR_S300 <= (others => '0');
		P_HR_S301 <= (others => '0');
		P_HR_S302 <= (others => '0');
		P_HR_S303 <= (others => '0');
		P_HR_S304 <= (others => '0');
		P_HR_S305 <= (others => '0');
		P_HR_S306 <= (others => '0');
		P_HR_S307 <= (others => '0');
		P_HR_S308 <= (others => '0');
		P_HR_S309 <= (others => '0');
		P_HR_S310 <= (others => '0');
		P_HR_S311 <= (others => '0');
		P_HR_S312 <= (others => '0');
		P_HR_S313 <= (others => '0');
		P_HR_S314 <= (others => '0');
		P_HR_S315 <= (others => '0');
		P_HR_S316 <= (others => '0');
		P_HR_S317 <= (others => '0');
		P_HR_S318 <= (others => '0');
		P_HR_S319 <= (others => '0');
		P_HR_S320 <= (others => '0');
		P_HR_S321 <= (others => '0');
		P_HR_S322 <= (others => '0');
		P_HR_S323 <= (others => '0');
		P_HR_S324 <= (others => '0');
		P_HR_S325 <= (others => '0');
		P_HR_S326 <= (others => '0');
		P_HR_S327 <= (others => '0');
		P_HR_S328 <= (others => '0');
		P_HR_S329 <= (others => '0');
		P_HR_S330 <= (others => '0');
		P_HR_S331 <= (others => '0');
		P_HR_S332 <= (others => '0');
		P_HR_S333 <= (others => '0');
		P_HR_S334 <= (others => '0');
		P_HR_S335 <= (others => '0');
		P_HR_S336 <= (others => '0');
		P_HR_S337 <= (others => '0');
		P_HR_S338 <= (others => '0');
		P_HR_S339 <= (others => '0');
		P_HR_S340 <= (others => '0');
		P_HR_S341 <= (others => '0');
		P_HR_S342 <= (others => '0');
		P_HR_S343 <= (others => '0');
		P_HR_S344 <= (others => '0');
		P_HR_S345 <= (others => '0');
		P_HR_S346 <= (others => '0');
		P_HR_S347 <= (others => '0');
		P_HR_S348 <= (others => '0');
		P_HR_S349 <= (others => '0');
		P_HR_S350 <= (others => '0');
		P_HR_S351 <= (others => '0');
		P_HR_S352 <= (others => '0');
		P_HR_S353 <= (others => '0');
		P_HR_S354 <= (others => '0');
		P_HR_S355 <= (others => '0');
		P_HR_S356 <= (others => '0');
		P_HR_S357 <= (others => '0');
		P_HR_S358 <= (others => '0');
		P_HR_S359 <= (others => '0');
		P_HR_S360 <= (others => '0');
		P_HR_S361 <= (others => '0');
		P_HR_S362 <= (others => '0');
		P_HR_S363 <= (others => '0');
		P_HR_S364 <= (others => '0');
		P_HR_S365 <= (others => '0');
		P_HR_S366 <= (others => '0');
		P_HR_S367 <= (others => '0');
		P_HR_S368 <= (others => '0');
		P_HR_S369 <= (others => '0');
		P_HR_S370 <= (others => '0');
		P_HR_S371 <= (others => '0');
		P_HR_S372 <= (others => '0');
		P_HR_S373 <= (others => '0');
		P_HR_S374 <= (others => '0');
		P_HR_S375 <= (others => '0');
		P_HR_S376 <= (others => '0');
		P_HR_S377 <= (others => '0');
		P_HR_S378 <= (others => '0');
		P_HR_S379 <= (others => '0');
		P_HR_S380 <= (others => '0');
		P_HR_S381 <= (others => '0');
		P_HR_S382 <= (others => '0');
		P_HR_S383 <= (others => '0');
		P_HR_S384 <= (others => '0');
		P_HR_S385 <= (others => '0');
		P_HR_S386 <= (others => '0');
		P_HR_S387 <= (others => '0');
		P_HR_S388 <= (others => '0');
		P_HR_S389 <= (others => '0');
		P_HR_S390 <= (others => '0');
		P_HR_S391 <= (others => '0');
		P_HR_S392 <= (others => '0');
		P_HR_S393 <= (others => '0');
		P_HR_S394 <= (others => '0');
		P_HR_S395 <= (others => '0');
		P_HR_S396 <= (others => '0');
		P_HR_S397 <= (others => '0');
		P_HR_S398 <= (others => '0');
		P_HR_S399 <= (others => '0');
		P_HR_S400 <= (others => '0');
		P_HR_S401 <= (others => '0');
		P_HR_S402 <= (others => '0');
		P_HR_S403 <= (others => '0');
		P_HR_S404 <= (others => '0');
		P_HR_S405 <= (others => '0');
		P_HR_S406 <= (others => '0');
		P_HR_S407 <= (others => '0');
		P_HR_S408 <= (others => '0');
		P_HR_S409 <= (others => '0');
		P_HR_S410 <= (others => '0');
		P_HR_S411 <= (others => '0');
		P_HR_S412 <= (others => '0');
		P_HR_S413 <= (others => '0');
		P_HR_S414 <= (others => '0');
		P_HR_S415 <= (others => '0');
		P_HR_S416 <= (others => '0');
		P_HR_S417 <= (others => '0');
		P_HR_S418 <= (others => '0');
		P_HR_S419 <= (others => '0');
		P_HR_S420 <= (others => '0');
		P_HR_S421 <= (others => '0');
		P_HR_S422 <= (others => '0');
		P_HR_S423 <= (others => '0');
		P_HR_S424 <= (others => '0');
		P_HR_S425 <= (others => '0');
		P_HR_S426 <= (others => '0');
		P_HR_S427 <= (others => '0');
		P_HR_S428 <= (others => '0');
			
		P_TEMP_S <= (others => '0');	
		P_EDA_S <= (others => '0');	
		P_HR_S <= (others => '0');		
	    
	    stress_score <= (others => '0');
			
		elsif (rising_edge(clk)) then
		
		if (state = NORMAL) then
		
			case temp is
				when "011110111" => P_TEMP_S <= "000000000010" + P_TEMP_S1;
				when "011111000" => P_TEMP_S <= "000110110110" + P_TEMP_S2;
				when "011111001" => P_TEMP_S <= "011001111011" + P_TEMP_S3;
				when "011111010" => P_TEMP_S <= "010111111010" + P_TEMP_S4;
				when "011111011" => P_TEMP_S <= "010011010100" + P_TEMP_S5;
				when "011111100" => P_TEMP_S <= "000000010111" + P_TEMP_S6;
				when "011111101" => P_TEMP_S <= "000000000010" + P_TEMP_S7;
				when "011111110" => P_TEMP_S <= "000110111001" + P_TEMP_S8;
				when "011111111" => P_TEMP_S <= "010010101101" + P_TEMP_S9;
				when "100000000" => P_TEMP_S <= "000111011010" + P_TEMP_S10;
				when "100000001" => P_TEMP_S <= "001000010011" + P_TEMP_S11;
				when "100000010" => P_TEMP_S <= "000101000100" + P_TEMP_S12;
				when "100000011" => P_TEMP_S <= "000010001000" + P_TEMP_S13;
				when "100000100" => P_TEMP_S <= "000001011111" + P_TEMP_S14;
				when "100000101" => P_TEMP_S <= "000001010101" + P_TEMP_S15;
				when "100000110" => P_TEMP_S <= "000001010000" + P_TEMP_S16;
				when "100000111" => P_TEMP_S <= "000001010011" + P_TEMP_S17;
				when "100001000" => P_TEMP_S <= "000001001101" + P_TEMP_S18;
				when "100001001" => P_TEMP_S <= "000001001000" + P_TEMP_S19;
				when "100001010" => P_TEMP_S <= "000001010010" + P_TEMP_S20;
				when "100001011" => P_TEMP_S <= "000011110111" + P_TEMP_S21;
				when "100001100" => P_TEMP_S <= "000100001101" + P_TEMP_S22;
				when "100001101" => P_TEMP_S <= "000100101011" + P_TEMP_S23;
				when "100001110" => P_TEMP_S <= "000010000001" + P_TEMP_S24;
				when "100001111" => P_TEMP_S <= "000010100011" + P_TEMP_S25;
				when "100010000" => P_TEMP_S <= "000000111000" + P_TEMP_S26;
				when "100010001" => P_TEMP_S <= "000000111101" + P_TEMP_S27;
				when "100010010" => P_TEMP_S <= "000001001110" + P_TEMP_S28;
				when "100010011" => P_TEMP_S <= "000010000000" + P_TEMP_S29;
				when "100010100" => P_TEMP_S <= "000000000010" + P_TEMP_S30;
				when others => P_TEMP_S      <= "000000000001";
			end case;
			
			
			case eda is
				when "0001000" => P_EDA_S <= "000000000010" + P_EDA_S1;
				when "0001001" => P_EDA_S <= "000101000011" + P_EDA_S2;
				when "0001010" => P_EDA_S <= "010001110100" + P_EDA_S3;
				when "0001011" => P_EDA_S <= "001000110001" + P_EDA_S4;
				when "0001100" => P_EDA_S <= "001010111100" + P_EDA_S5;
				when "0001101" => P_EDA_S <= "000001011111" + P_EDA_S6;
				when "0001110" => P_EDA_S <= "000100000110" + P_EDA_S7;
				when "0001111" => P_EDA_S <= "000101001010" + P_EDA_S8;
				when "0010000" => P_EDA_S <= "000001010111" + P_EDA_S9;
				when "0010001" => P_EDA_S <= "000000000101" + P_EDA_S10;
				when "0010010" => P_EDA_S <= "000001111011" + P_EDA_S11;
				when "0010011" => P_EDA_S <= "000010011101" + P_EDA_S12;
				when "0010100" => P_EDA_S <= "000010000101" + P_EDA_S13;
				when "0010101" => P_EDA_S <= "000100100011" + P_EDA_S14;
				when "0010110" => P_EDA_S <= "000010001010" + P_EDA_S15;
				when "0010111" => P_EDA_S <= "000100010100" + P_EDA_S16;
				when "0011000" => P_EDA_S <= "000010011001" + P_EDA_S17;
				when "0011001" => P_EDA_S <= "000001001100" + P_EDA_S18;
				when "0011010" => P_EDA_S <= "000000010011" + P_EDA_S19;
				when "0011011" => P_EDA_S <= "000000001111" + P_EDA_S20;
				when "0011100" => P_EDA_S <= "000000000001" + P_EDA_S21;
				when "0110110" => P_EDA_S <= "000000000010" + P_EDA_S22;
				when "0110111" => P_EDA_S <= "000100100111" + P_EDA_S23;
				when "0111000" => P_EDA_S <= "000010101100" + P_EDA_S24;
				when "0111001" => P_EDA_S <= "000000011001" + P_EDA_S25;
				when "0111010" => P_EDA_S <= "000001100010" + P_EDA_S26;
				when "0111011" => P_EDA_S <= "000010101101" + P_EDA_S27;
				when "0111100" => P_EDA_S <= "000100001100" + P_EDA_S28;
				when "0111101" => P_EDA_S <= "000010111100" + P_EDA_S29;
				when "0111110" => P_EDA_S <= "000101110000" + P_EDA_S30;
				when "0111111" => P_EDA_S <= "000110100010" + P_EDA_S31;
				when "1000000" => P_EDA_S <= "000100000100" + P_EDA_S32;
				when "1000001" => P_EDA_S <= "000101100100" + P_EDA_S33;
				when "1000010" => P_EDA_S <= "000101000000" + P_EDA_S34;
				when "1000011" => P_EDA_S <= "000100001101" + P_EDA_S35;
				when "1000100" => P_EDA_S <= "000011111111" + P_EDA_S36;
				when "1000101" => P_EDA_S <= "000001111100" + P_EDA_S37;
				when "1000110" => P_EDA_S <= "000010101110" + P_EDA_S38;
				when "1000111" => P_EDA_S <= "000001101001" + P_EDA_S39;
				when "1001000" => P_EDA_S <= "000001101111" + P_EDA_S40;
				when "1001001" => P_EDA_S <= "000001010110" + P_EDA_S41;
				when "1001010" => P_EDA_S <= "000001110111" + P_EDA_S42;
				when "1001011" => P_EDA_S <= "000001111111" + P_EDA_S43;
				when "1001100" => P_EDA_S <= "000101001010" + P_EDA_S44;
				when "1001101" => P_EDA_S <= "000001101000" + P_EDA_S45;
				when "1001110" => P_EDA_S <= "000000000110" + P_EDA_S46;
				when "1001111" => P_EDA_S <= "000000000101" + P_EDA_S47;
				when "1010000" => P_EDA_S <= "000000000101" + P_EDA_S48;
				when "1010001" => P_EDA_S <= "000000001100" + P_EDA_S49;
				when "1010010" => P_EDA_S <= "000000010011" + P_EDA_S50;
				when "1010011" => P_EDA_S <= "000000001110" + P_EDA_S51;
				when "1010100" => P_EDA_S <= "000000001111" + P_EDA_S52;
				when "1010101" => P_EDA_S <= "000000100000" + P_EDA_S53;
				when "1010110" => P_EDA_S <= "000000100111" + P_EDA_S54;
				when "1010111" => P_EDA_S <= "000000100001" + P_EDA_S55;
				when "1011000" => P_EDA_S <= "000000011110" + P_EDA_S56;
				when "1011001" => P_EDA_S <= "000000001111" + P_EDA_S57;
				when "1011010" => P_EDA_S <= "000000010100" + P_EDA_S58;
				when "1011011" => P_EDA_S <= "000000011110" + P_EDA_S59;
				when "1011100" => P_EDA_S <= "000000001110" + P_EDA_S60;
				when "1011101" => P_EDA_S <= "000000001001" + P_EDA_S61;
				when "1011110" => P_EDA_S <= "000000001101" + P_EDA_S62;
				when "1011111" => P_EDA_S <= "000000100011" + P_EDA_S63;
				when "1100000" => P_EDA_S <= "000000010010" + P_EDA_S64;
				when "1100001" => P_EDA_S <= "000000000010" + P_EDA_S65;
				when others    => P_EDA_S <= "000000000001";
			end case;

			case hr is
				when "00000001100" => P_HR_S <= "000000001001" + P_HR_S1;
				when "00000001110" => P_HR_S <= "000000001001" + P_HR_S2;
				when "00000010011" => P_HR_S <= "000000001001" + P_HR_S3;
				when "00000010111" => P_HR_S <= "000000001001" + P_HR_S4;
				when "00000011001" => P_HR_S <= "000000001001" + P_HR_S5;
				when "00000011100" => P_HR_S <= "000000001001" + P_HR_S6;
				when "00000100101" => P_HR_S <= "000000001001" + P_HR_S7;
				when "00000100110" => P_HR_S <= "000000001001" + P_HR_S8;
				when "00000110001" => P_HR_S <= "000000001001" + P_HR_S9;
				when "00001000111" => P_HR_S <= "000000001001" + P_HR_S10;
				when "00001001100" => P_HR_S <= "000000001001" + P_HR_S11;
				when "00001001101" => P_HR_S <= "000000001001" + P_HR_S12;
				when "00001001110" => P_HR_S <= "000000001001" + P_HR_S13;
				when "00001010001" => P_HR_S <= "000000001001" + P_HR_S14;
				when "00001010101" => P_HR_S <= "000000010010" + P_HR_S15;
				when "00001010111" => P_HR_S <= "000000001001" + P_HR_S16;
				when "00001011001" => P_HR_S <= "000000010010" + P_HR_S17;
				when "00001100001" => P_HR_S <= "000000001001" + P_HR_S18;
				when "00001100010" => P_HR_S <= "000000001001" + P_HR_S19;
				when "00001100011" => P_HR_S <= "000000001001" + P_HR_S20;
				when "00001110000" => P_HR_S <= "000000001001" + P_HR_S21;
				when "00001110001" => P_HR_S <= "000000001001" + P_HR_S22;
				when "00001110101" => P_HR_S <= "000000001001" + P_HR_S23;
				when "00001111000" => P_HR_S <= "000000001001" + P_HR_S24;
				when "00001111100" => P_HR_S <= "000000001001" + P_HR_S25;
				when "00001111111" => P_HR_S <= "000000100011" + P_HR_S26;
				when "00010000011" => P_HR_S <= "000000001001" + P_HR_S27;
				when "00010000111" => P_HR_S <= "000000001001" + P_HR_S28;
				when "00010001011" => P_HR_S <= "000000001001" + P_HR_S29;
				when "00010001110" => P_HR_S <= "000000001001" + P_HR_S30;
				when "00010001111" => P_HR_S <= "000000001001" + P_HR_S31;
				when "00010010000" => P_HR_S <= "000000010010" + P_HR_S32;
				when "00010010010" => P_HR_S <= "000000001001" + P_HR_S33;
				when "00010010011" => P_HR_S <= "000000001001" + P_HR_S34;
				when "00010010100" => P_HR_S <= "000000001001" + P_HR_S35;
				when "00010010101" => P_HR_S <= "000000001001" + P_HR_S36;
				when "00010011000" => P_HR_S <= "000000001001" + P_HR_S37;
				when "00010011110" => P_HR_S <= "000000001001" + P_HR_S38;
				when "00010100010" => P_HR_S <= "000000001001" + P_HR_S39;
				when "00010110101" => P_HR_S <= "000000001001" + P_HR_S40;
				when "00010110110" => P_HR_S <= "000000010010" + P_HR_S41;
				when "00010111000" => P_HR_S <= "000000001001" + P_HR_S42;
				when "00010111001" => P_HR_S <= "000000001001" + P_HR_S43;
				when "00010111100" => P_HR_S <= "000000001001" + P_HR_S44;
				when "00010111101" => P_HR_S <= "000000001001" + P_HR_S45;
				when "00010111110" => P_HR_S <= "000000001001" + P_HR_S46;
				when "00010111111" => P_HR_S <= "000000001001" + P_HR_S47;
				when "00011000000" => P_HR_S <= "000000010010" + P_HR_S48;
				when "00011000001" => P_HR_S <= "000000001001" + P_HR_S49;
				when "00011000101" => P_HR_S <= "000000010010" + P_HR_S50;
				when "00011000110" => P_HR_S <= "000000010010" + P_HR_S51;
				when "00011000111" => P_HR_S <= "000000001001" + P_HR_S52;
				when "00011001000" => P_HR_S <= "000000001001" + P_HR_S53;
				when "00011001001" => P_HR_S <= "000000001001" + P_HR_S54;
				when "00011001010" => P_HR_S <= "000000011010" + P_HR_S55;
				when "00011001011" => P_HR_S <= "000000010010" + P_HR_S56;
				when "00011001101" => P_HR_S <= "000000010010" + P_HR_S57;
				when "00011001110" => P_HR_S <= "000000010010" + P_HR_S58;
				when "00011010000" => P_HR_S <= "000000010010" + P_HR_S59;
				when "00011010001" => P_HR_S <= "000000010010" + P_HR_S60;
				when "00011010100" => P_HR_S <= "000000001001" + P_HR_S61;
				when "00011011010" => P_HR_S <= "000000001001" + P_HR_S62;
				when "00011100100" => P_HR_S <= "000000001001" + P_HR_S63;
				when "00011111001" => P_HR_S <= "000000001001" + P_HR_S64;
				when "00100001111" => P_HR_S <= "000000001001" + P_HR_S65;
				when "00100010000" => P_HR_S <= "000000011010" + P_HR_S66;
				when "00100010001" => P_HR_S <= "000000001001" + P_HR_S67;
				when "00100010100" => P_HR_S <= "000000001001" + P_HR_S68;
				when "00100011001" => P_HR_S <= "000000001001" + P_HR_S69;
				when "00100011011" => P_HR_S <= "000000001001" + P_HR_S70;
				when "00100011100" => P_HR_S <= "000000001001" + P_HR_S71;
				when "00100011110" => P_HR_S <= "000000001001" + P_HR_S72;
				when "00100011111" => P_HR_S <= "000000001001" + P_HR_S73;
				when "00100100000" => P_HR_S <= "000000100011" + P_HR_S74;
				when "00100100001" => P_HR_S <= "000000001001" + P_HR_S75;
				when "00100100010" => P_HR_S <= "000000001001" + P_HR_S76;
				when "00100100011" => P_HR_S <= "000000001001" + P_HR_S77;
				when "00100100100" => P_HR_S <= "000000001001" + P_HR_S78;
				when "00100100101" => P_HR_S <= "000000001001" + P_HR_S79;
				when "00100100110" => P_HR_S <= "000000001001" + P_HR_S80;
				when "00100100111" => P_HR_S <= "000000001001" + P_HR_S81;
				when "00100101010" => P_HR_S <= "000000001001" + P_HR_S82;
				when "00100101100" => P_HR_S <= "000000010010" + P_HR_S83;
				when "00100101110" => P_HR_S <= "000000001001" + P_HR_S84;
				when "00100110010" => P_HR_S <= "000000001001" + P_HR_S85;
				when "00100110011" => P_HR_S <= "000000001001" + P_HR_S86;
				when "00100110100" => P_HR_S <= "000000001001" + P_HR_S87;
				when "00100110111" => P_HR_S <= "000000010010" + P_HR_S88;
				when "00100111000" => P_HR_S <= "000000001001" + P_HR_S89;
				when "00100111001" => P_HR_S <= "000000001001" + P_HR_S90;
				when "00100111101" => P_HR_S <= "000000010010" + P_HR_S91;
				when "00101000101" => P_HR_S <= "000000001001" + P_HR_S92;
				when "00101001101" => P_HR_S <= "000000001001" + P_HR_S93;
				when "00101010010" => P_HR_S <= "000000001001" + P_HR_S94;
				when "00101010100" => P_HR_S <= "000000001001" + P_HR_S95;
				when "00101011001" => P_HR_S <= "000000001001" + P_HR_S96;
				when "00110010011" => P_HR_S <= "000000001001" + P_HR_S97;
				when "00110010111" => P_HR_S <= "000000001001" + P_HR_S98;
				when "00110011000" => P_HR_S <= "000000001001" + P_HR_S99;
				when "00110011001" => P_HR_S <= "000000001001" + P_HR_S100;
				when "00110110011" => P_HR_S <= "000000010010" + P_HR_S101;
				when "00110110110" => P_HR_S <= "000000001001" + P_HR_S102;
				when "00110111100" => P_HR_S <= "000000010010" + P_HR_S103;
				when "00110111110" => P_HR_S <= "000000001001" + P_HR_S104;
				when "00111000000" => P_HR_S <= "000000001001" + P_HR_S105;
				when "00111000010" => P_HR_S <= "000000001001" + P_HR_S106;
				when "00111000011" => P_HR_S <= "000000001001" + P_HR_S107;
				when "00111000111" => P_HR_S <= "000000010010" + P_HR_S108;
				when "00111001001" => P_HR_S <= "000000010010" + P_HR_S109;
				when "00111001100" => P_HR_S <= "000000001001" + P_HR_S110;
				when "00111001101" => P_HR_S <= "000000001001" + P_HR_S111;
				when "00111001111" => P_HR_S <= "000000001001" + P_HR_S112;
				when "00111010010" => P_HR_S <= "000000001001" + P_HR_S113;
				when "00111010101" => P_HR_S <= "000000001001" + P_HR_S114;
				when "00111010111" => P_HR_S <= "000000001001" + P_HR_S115;
				when "00111011000" => P_HR_S <= "000000001001" + P_HR_S116;
				when "00111011001" => P_HR_S <= "000000001001" + P_HR_S117;
				when "00111011100" => P_HR_S <= "000000011010" + P_HR_S118;
				when "00111011101" => P_HR_S <= "000000011010" + P_HR_S119;
				when "00111100001" => P_HR_S <= "000000011010" + P_HR_S120;
				when "00111100011" => P_HR_S <= "000000001001" + P_HR_S121;
				when "00111100110" => P_HR_S <= "000000001001" + P_HR_S122;
				when "00111101011" => P_HR_S <= "000000001001" + P_HR_S123;
				when "00111101111" => P_HR_S <= "000000010010" + P_HR_S124;
				when "00111110000" => P_HR_S <= "000000001001" + P_HR_S125;
				when "00111110010" => P_HR_S <= "000000001001" + P_HR_S126;
				when "00111110100" => P_HR_S <= "000000001001" + P_HR_S127;
				when "00111110101" => P_HR_S <= "000000010010" + P_HR_S128;
				when "00111110110" => P_HR_S <= "000000011010" + P_HR_S129;
				when "00111111000" => P_HR_S <= "000000001001" + P_HR_S130;
				when "00111111001" => P_HR_S <= "000000010010" + P_HR_S131;
				when "00111111100" => P_HR_S <= "000000011010" + P_HR_S132;
				when "00111111111" => P_HR_S <= "000000001001" + P_HR_S133;
				when "01000000011" => P_HR_S <= "000000010010" + P_HR_S134;
				when "01000000100" => P_HR_S <= "000000010010" + P_HR_S135;
				when "01000000101" => P_HR_S <= "000000001001" + P_HR_S136;
				when "01000000110" => P_HR_S <= "000000010010" + P_HR_S137;
				when "01000000111" => P_HR_S <= "000000010010" + P_HR_S138;
				when "01000001001" => P_HR_S <= "000000001001" + P_HR_S139;
				when "01000001010" => P_HR_S <= "000000001001" + P_HR_S140;
				when "01000001011" => P_HR_S <= "000000001001" + P_HR_S141;
				when "01000001101" => P_HR_S <= "000000001001" + P_HR_S142;
				when "01000001111" => P_HR_S <= "000000101100" + P_HR_S143;
				when "01000010001" => P_HR_S <= "000000100011" + P_HR_S144;
				when "01000010010" => P_HR_S <= "000000010010" + P_HR_S145;
				when "01000010100" => P_HR_S <= "000000110101" + P_HR_S146;
				when "01000010101" => P_HR_S <= "000000001001" + P_HR_S147;
				when "01000010110" => P_HR_S <= "000000011010" + P_HR_S148;
				when "01000010111" => P_HR_S <= "000000001001" + P_HR_S149;
				when "01000011000" => P_HR_S <= "000000001001" + P_HR_S150;
				when "01000011010" => P_HR_S <= "000000100011" + P_HR_S151;
				when "01000011011" => P_HR_S <= "000000011010" + P_HR_S152;
				when "01000011100" => P_HR_S <= "000000001001" + P_HR_S153;
				when "01000011101" => P_HR_S <= "000000100011" + P_HR_S154;
				when "01000011111" => P_HR_S <= "000000001001" + P_HR_S155;
				when "01000100000" => P_HR_S <= "000000010010" + P_HR_S156;
				when "01000100001" => P_HR_S <= "000000011010" + P_HR_S157;
				when "01000100011" => P_HR_S <= "000000001001" + P_HR_S158;
				when "01000100100" => P_HR_S <= "000000001001" + P_HR_S159;
				when "01000100111" => P_HR_S <= "000000001001" + P_HR_S160;
				when "01000101000" => P_HR_S <= "000000010010" + P_HR_S161;
				when "01000101001" => P_HR_S <= "000000001001" + P_HR_S162;
				when "01000101010" => P_HR_S <= "000000101100" + P_HR_S163;
				when "01000101011" => P_HR_S <= "000000101100" + P_HR_S164;
				when "01000101100" => P_HR_S <= "000000011010" + P_HR_S165;
				when "01000101101" => P_HR_S <= "000000010010" + P_HR_S166;
				when "01000101110" => P_HR_S <= "000000011010" + P_HR_S167;
				when "01000101111" => P_HR_S <= "000000101100" + P_HR_S168;
				when "01000110000" => P_HR_S <= "000000001001" + P_HR_S169;
				when "01000110001" => P_HR_S <= "000000010010" + P_HR_S170;
				when "01000110011" => P_HR_S <= "000000101100" + P_HR_S171;
				when "01000110100" => P_HR_S <= "000000001001" + P_HR_S172;
				when "01000110101" => P_HR_S <= "000000001001" + P_HR_S173;
				when "01000110110" => P_HR_S <= "000000011010" + P_HR_S174;
				when "01000110111" => P_HR_S <= "000000001001" + P_HR_S175;
				when "01000111000" => P_HR_S <= "000000010010" + P_HR_S176;
				when "01000111001" => P_HR_S <= "000001100001" + P_HR_S177;
				when "01000111010" => P_HR_S <= "000000101100" + P_HR_S178;
				when "01000111011" => P_HR_S <= "000000001001" + P_HR_S179;
				when "01000111100" => P_HR_S <= "000000001001" + P_HR_S180;
				when "01000111101" => P_HR_S <= "000000101100" + P_HR_S181;
				when "01000111110" => P_HR_S <= "000000100011" + P_HR_S182;
				when "01000111111" => P_HR_S <= "000000010010" + P_HR_S183;
				when "01001000000" => P_HR_S <= "000000100011" + P_HR_S184;
				when "01001000001" => P_HR_S <= "000000011010" + P_HR_S185;
				when "01001000010" => P_HR_S <= "000000111110" + P_HR_S186;
				when "01001000011" => P_HR_S <= "000000011010" + P_HR_S187;
				when "01001000100" => P_HR_S <= "000000111110" + P_HR_S188;
				when "01001000101" => P_HR_S <= "000000011010" + P_HR_S189;
				when "01001000110" => P_HR_S <= "000000011010" + P_HR_S190;
				when "01001000111" => P_HR_S <= "000000011010" + P_HR_S191;
				when "01001001000" => P_HR_S <= "000000001001" + P_HR_S192;
				when "01001001001" => P_HR_S <= "000000011010" + P_HR_S193;
				when "01001001010" => P_HR_S <= "000000010010" + P_HR_S194;
				when "01001001011" => P_HR_S <= "000000011010" + P_HR_S195;
				when "01001001100" => P_HR_S <= "000000011010" + P_HR_S196;
				when "01001001101" => P_HR_S <= "000000110101" + P_HR_S197;
				when "01001001111" => P_HR_S <= "000000001001" + P_HR_S198;
				when "01001010001" => P_HR_S <= "000000010010" + P_HR_S199;
				when "01001010010" => P_HR_S <= "000000011010" + P_HR_S200;
				when "01001010011" => P_HR_S <= "000000001001" + P_HR_S201;
				when "01001010100" => P_HR_S <= "000000111110" + P_HR_S202;
				when "01001010101" => P_HR_S <= "000000001001" + P_HR_S203;
				when "01001010110" => P_HR_S <= "000000011010" + P_HR_S204;
				when "01001010111" => P_HR_S <= "000000001001" + P_HR_S205;
				when "01001011000" => P_HR_S <= "000000001001" + P_HR_S206;
				when "01001011001" => P_HR_S <= "000000001001" + P_HR_S207;
				when "01001011010" => P_HR_S <= "000000101100" + P_HR_S208;
				when "01001011011" => P_HR_S <= "000000011010" + P_HR_S209;
				when "01001011100" => P_HR_S <= "000000001001" + P_HR_S210;
				when "01001011101" => P_HR_S <= "000000110101" + P_HR_S211;
				when "01001011110" => P_HR_S <= "000000101100" + P_HR_S212;
				when "01001100001" => P_HR_S <= "000000010010" + P_HR_S213;
				when "01001100010" => P_HR_S <= "000000011010" + P_HR_S214;
				when "01001100011" => P_HR_S <= "000000011010" + P_HR_S215;
				when "01001100100" => P_HR_S <= "000000010010" + P_HR_S216;
				when "01001100101" => P_HR_S <= "000000101100" + P_HR_S217;
				when "01001100110" => P_HR_S <= "000000100011" + P_HR_S218;
				when "01001100111" => P_HR_S <= "000000010010" + P_HR_S219;
				when "01001101001" => P_HR_S <= "000000001001" + P_HR_S220;
				when "01001101010" => P_HR_S <= "000000001001" + P_HR_S221;
				when "01001101011" => P_HR_S <= "000000101100" + P_HR_S222;
				when "01001101100" => P_HR_S <= "000000101100" + P_HR_S223;
				when "01001101101" => P_HR_S <= "000000011010" + P_HR_S224;
				when "01001101110" => P_HR_S <= "000000011010" + P_HR_S225;
				when "01001101111" => P_HR_S <= "000000001001" + P_HR_S226;
				when "01001110001" => P_HR_S <= "000000100011" + P_HR_S227;
				when "01001110011" => P_HR_S <= "000000010010" + P_HR_S228;
				when "01001110100" => P_HR_S <= "000000010010" + P_HR_S229;
				when "01001110101" => P_HR_S <= "000000011010" + P_HR_S230;
				when "01001110110" => P_HR_S <= "000000100011" + P_HR_S231;
				when "01001111000" => P_HR_S <= "000000010010" + P_HR_S232;
				when "01001111001" => P_HR_S <= "000000011010" + P_HR_S233;
				when "01001111010" => P_HR_S <= "000000100011" + P_HR_S234;
				when "01001111011" => P_HR_S <= "000000011010" + P_HR_S235;
				when "01001111100" => P_HR_S <= "000000001001" + P_HR_S236;
				when "01001111110" => P_HR_S <= "000001001111" + P_HR_S237;
				when "01001111111" => P_HR_S <= "000000100011" + P_HR_S238;
				when "01010000000" => P_HR_S <= "000000110101" + P_HR_S239;
				when "01010000001" => P_HR_S <= "000000101100" + P_HR_S240;
				when "01010000010" => P_HR_S <= "000000110101" + P_HR_S241;
				when "01010000100" => P_HR_S <= "000000011010" + P_HR_S242;
				when "01010000101" => P_HR_S <= "000000101100" + P_HR_S243;
				when "01010000110" => P_HR_S <= "000000101100" + P_HR_S244;
				when "01010001001" => P_HR_S <= "000000101100" + P_HR_S245;
				when "01010001010" => P_HR_S <= "000000011010" + P_HR_S246;
				when "01010001011" => P_HR_S <= "000000010010" + P_HR_S247;
				when "01010001110" => P_HR_S <= "000000011010" + P_HR_S248;
				when "01010001111" => P_HR_S <= "000000111110" + P_HR_S249;
				when "01010010000" => P_HR_S <= "000000001001" + P_HR_S250;
				when "01010010010" => P_HR_S <= "000001000110" + P_HR_S251;
				when "01010010011" => P_HR_S <= "000000010010" + P_HR_S252;
				when "01010010100" => P_HR_S <= "000000010010" + P_HR_S253;
				when "01010010101" => P_HR_S <= "000000010010" + P_HR_S254;
				when "01010010111" => P_HR_S <= "000000001001" + P_HR_S255;
				when "01010011000" => P_HR_S <= "000000011010" + P_HR_S256;
				when "01010011001" => P_HR_S <= "000000011010" + P_HR_S257;
				when "01010011011" => P_HR_S <= "000000101100" + P_HR_S258;
				when "01010011100" => P_HR_S <= "000000110101" + P_HR_S259;
				when "01010011101" => P_HR_S <= "000000010010" + P_HR_S260;
				when "01010011111" => P_HR_S <= "000000100011" + P_HR_S261;
				when "01010100000" => P_HR_S <= "000000110101" + P_HR_S262;
				when "01010100001" => P_HR_S <= "000000011010" + P_HR_S263;
				when "01010100011" => P_HR_S <= "000000011010" + P_HR_S264;
				when "01010100100" => P_HR_S <= "000000010010" + P_HR_S265;
				when "01010100101" => P_HR_S <= "000000001001" + P_HR_S266;
				when "01010100111" => P_HR_S <= "000001001111" + P_HR_S267;
				when "01010101000" => P_HR_S <= "000000010010" + P_HR_S268;
				when "01010101010" => P_HR_S <= "000000010010" + P_HR_S269;
				when "01010101011" => P_HR_S <= "000000010010" + P_HR_S270;
				when "01010101100" => P_HR_S <= "000000110101" + P_HR_S271;
				when "01010101110" => P_HR_S <= "000000101100" + P_HR_S272;
				when "01010101111" => P_HR_S <= "000000011010" + P_HR_S273;
				when "01010110001" => P_HR_S <= "000000010010" + P_HR_S274;
				when "01010110010" => P_HR_S <= "000000011010" + P_HR_S275;
				when "01010110011" => P_HR_S <= "000000010010" + P_HR_S276;
				when "01010110101" => P_HR_S <= "000000011010" + P_HR_S277;
				when "01010110110" => P_HR_S <= "000000100011" + P_HR_S278;
				when "01010111000" => P_HR_S <= "000000010010" + P_HR_S279;
				when "01010111001" => P_HR_S <= "000000110101" + P_HR_S280;
				when "01010111100" => P_HR_S <= "000000111110" + P_HR_S281;
				when "01010111101" => P_HR_S <= "000000011010" + P_HR_S282;
				when "01010111111" => P_HR_S <= "000000101100" + P_HR_S283;
				when "01011000000" => P_HR_S <= "000000010010" + P_HR_S284;
				when "01011000010" => P_HR_S <= "000000010010" + P_HR_S285;
				when "01011000011" => P_HR_S <= "000000011010" + P_HR_S286;
				when "01011000101" => P_HR_S <= "000000111110" + P_HR_S287;
				when "01011000110" => P_HR_S <= "000000100011" + P_HR_S288;
				when "01011001000" => P_HR_S <= "000000100011" + P_HR_S289;
				when "01011001001" => P_HR_S <= "000000010010" + P_HR_S290;
				when "01011001011" => P_HR_S <= "000000010010" + P_HR_S291;
				when "01011001100" => P_HR_S <= "000000011010" + P_HR_S292;
				when "01011001110" => P_HR_S <= "000001000110" + P_HR_S293;
				when "01011001111" => P_HR_S <= "000000101100" + P_HR_S294;
				when "01011010001" => P_HR_S <= "000000110101" + P_HR_S295;
				when "01011010011" => P_HR_S <= "000000010010" + P_HR_S296;
				when "01011010100" => P_HR_S <= "000000100011" + P_HR_S297;
				when "01011010110" => P_HR_S <= "000000111110" + P_HR_S298;
				when "01011010111" => P_HR_S <= "000000100011" + P_HR_S299;
				when "01011011001" => P_HR_S <= "000000110101" + P_HR_S300;
				when "01011011010" => P_HR_S <= "000000100011" + P_HR_S301;
				when "01011011100" => P_HR_S <= "000000010010" + P_HR_S302;
				when "01011011110" => P_HR_S <= "000000101100" + P_HR_S303;
				when "01011011111" => P_HR_S <= "000000110101" + P_HR_S304;
				when "01011100001" => P_HR_S <= "000000101100" + P_HR_S305;
				when "01011100010" => P_HR_S <= "000000011010" + P_HR_S306;
				when "01011100100" => P_HR_S <= "000000011010" + P_HR_S307;
				when "01011100110" => P_HR_S <= "000000100011" + P_HR_S308;
				when "01011100111" => P_HR_S <= "000001000110" + P_HR_S309;
				when "01011101001" => P_HR_S <= "000000110101" + P_HR_S310;
				when "01011101011" => P_HR_S <= "000000100011" + P_HR_S311;
				when "01011101100" => P_HR_S <= "000000110101" + P_HR_S312;
				when "01011101110" => P_HR_S <= "000000111110" + P_HR_S313;
				when "01011110000" => P_HR_S <= "000000110101" + P_HR_S314;
				when "01011110001" => P_HR_S <= "000000001001" + P_HR_S315;
				when "01011110011" => P_HR_S <= "000000011010" + P_HR_S316;
				when "01011110101" => P_HR_S <= "000000110101" + P_HR_S317;
				when "01011110110" => P_HR_S <= "000000110101" + P_HR_S318;
				when "01011111000" => P_HR_S <= "000000011010" + P_HR_S319;
				when "01011111010" => P_HR_S <= "000000101100" + P_HR_S320;
				when "01011111100" => P_HR_S <= "000000110101" + P_HR_S321;
				when "01011111101" => P_HR_S <= "000001101001" + P_HR_S322;
				when "01011111111" => P_HR_S <= "000000010010" + P_HR_S323;
				when "01100000001" => P_HR_S <= "000000100011" + P_HR_S324;
				when "01100000011" => P_HR_S <= "000000001001" + P_HR_S325;
				when "01100000100" => P_HR_S <= "000000111110" + P_HR_S326;
				when "01100000110" => P_HR_S <= "000000100011" + P_HR_S327;
				when "01100001000" => P_HR_S <= "000001001111" + P_HR_S328;
				when "01100001010" => P_HR_S <= "000000010010" + P_HR_S329;
				when "01100001100" => P_HR_S <= "000000100011" + P_HR_S330;
				when "01100001101" => P_HR_S <= "000000101100" + P_HR_S331;
				when "01100001111" => P_HR_S <= "000001000110" + P_HR_S332;
				when "01100010001" => P_HR_S <= "000000011010" + P_HR_S333;
				when "01100010011" => P_HR_S <= "000001000110" + P_HR_S334;
				when "01100010101" => P_HR_S <= "000000110101" + P_HR_S335;
				when "01100010111" => P_HR_S <= "000000011010" + P_HR_S336;
				when "01100011000" => P_HR_S <= "000000101100" + P_HR_S337;
				when "01100011010" => P_HR_S <= "000000111110" + P_HR_S338;
				when "01100011110" => P_HR_S <= "000000111110" + P_HR_S339;
				when "01100100000" => P_HR_S <= "000001001111" + P_HR_S340;
				when "01100100010" => P_HR_S <= "000000010010" + P_HR_S341;
				when "01100100100" => P_HR_S <= "000000001001" + P_HR_S342;
				when "01100100110" => P_HR_S <= "000000011010" + P_HR_S343;
				when "01100101000" => P_HR_S <= "000001011000" + P_HR_S344;
				when "01100101010" => P_HR_S <= "000001001111" + P_HR_S345;
				when "01100101100" => P_HR_S <= "000000011010" + P_HR_S346;
				when "01100101110" => P_HR_S <= "000000001001" + P_HR_S347;
				when "01100110000" => P_HR_S <= "000000010010" + P_HR_S348;
				when "01100110010" => P_HR_S <= "000000110101" + P_HR_S349;
				when "01100110100" => P_HR_S <= "000000011010" + P_HR_S350;
				when "01100110110" => P_HR_S <= "000000100011" + P_HR_S351;
				when "01100111000" => P_HR_S <= "000000011010" + P_HR_S352;
				when "01100111010" => P_HR_S <= "000000101100" + P_HR_S353;
				when "01100111100" => P_HR_S <= "000000011010" + P_HR_S354;
				when "01100111110" => P_HR_S <= "000000101100" + P_HR_S355;
				when "01101000000" => P_HR_S <= "000000110101" + P_HR_S356;
				when "01101000010" => P_HR_S <= "000000100011" + P_HR_S357;
				when "01101000100" => P_HR_S <= "000000100011" + P_HR_S358;
				when "01101000110" => P_HR_S <= "000000001001" + P_HR_S359;
				when "01101001000" => P_HR_S <= "000000010010" + P_HR_S360;
				when "01101001100" => P_HR_S <= "000000011010" + P_HR_S361;
				when "01101001110" => P_HR_S <= "000000101100" + P_HR_S362;
				when "01101010000" => P_HR_S <= "000000001001" + P_HR_S363;
				when "01101010011" => P_HR_S <= "000000101100" + P_HR_S364;
				when "01101010101" => P_HR_S <= "000000010010" + P_HR_S365;
				when "01101010111" => P_HR_S <= "000000001001" + P_HR_S366;
				when "01101011001" => P_HR_S <= "000000001001" + P_HR_S367;
				when "01101011011" => P_HR_S <= "000000100011" + P_HR_S368;
				when "01101011110" => P_HR_S <= "000000001001" + P_HR_S369;
				when "01101100000" => P_HR_S <= "000000011010" + P_HR_S370;
				when "01101100010" => P_HR_S <= "000000001001" + P_HR_S371;
				when "01101100100" => P_HR_S <= "000000100011" + P_HR_S372;
				when "01101100110" => P_HR_S <= "000000110101" + P_HR_S373;
				when "01101101001" => P_HR_S <= "000000011010" + P_HR_S374;
				when "01101101011" => P_HR_S <= "000000001001" + P_HR_S375;
				when "01101101101" => P_HR_S <= "000000010010" + P_HR_S376;
				when "01101110000" => P_HR_S <= "000000001001" + P_HR_S377;
				when "01101110010" => P_HR_S <= "000000010010" + P_HR_S378;
				when "01101110100" => P_HR_S <= "000000010010" + P_HR_S379;
				when "01101111011" => P_HR_S <= "000000010010" + P_HR_S380;
				when "01101111110" => P_HR_S <= "000000001001" + P_HR_S381;
				when "01110000101" => P_HR_S <= "000000001001" + P_HR_S382;
				when "01110000111" => P_HR_S <= "000000010010" + P_HR_S383;
				when "01110001010" => P_HR_S <= "000000010010" + P_HR_S384;
				when "01110001100" => P_HR_S <= "000000010010" + P_HR_S385;
				when "01110001111" => P_HR_S <= "000000010010" + P_HR_S386;
				when "01110010100" => P_HR_S <= "000000010010" + P_HR_S387;
				when "01110010110" => P_HR_S <= "000000001001" + P_HR_S388;
				when "01110011001" => P_HR_S <= "000000001001" + P_HR_S389;
				when "01110011011" => P_HR_S <= "000000001001" + P_HR_S390;
				when "01110100011" => P_HR_S <= "000000001001" + P_HR_S391;
				when "01110101101" => P_HR_S <= "000000001001" + P_HR_S392;
				when "01110110010" => P_HR_S <= "000000010010" + P_HR_S393;
				when "01110110101" => P_HR_S <= "000000001001" + P_HR_S394;
				when "01110111000" => P_HR_S <= "000000011010" + P_HR_S395;
				when "01110111011" => P_HR_S <= "000000001001" + P_HR_S396;
				when "01111000000" => P_HR_S <= "000000001001" + P_HR_S397;
				when "01111000110" => P_HR_S <= "000000001001" + P_HR_S398;
				when "01111001000" => P_HR_S <= "000000001001" + P_HR_S399;
				when "01111001011" => P_HR_S <= "000000010010" + P_HR_S400;
				when "01111001110" => P_HR_S <= "000000010010" + P_HR_S401;
				when "01111010001" => P_HR_S <= "000000010010" + P_HR_S402;
				when "01111010100" => P_HR_S <= "000000010010" + P_HR_S403;
				when "01111010110" => P_HR_S <= "000000001001" + P_HR_S404;
				when "01111011100" => P_HR_S <= "000000001001" + P_HR_S405;
				when "01111011111" => P_HR_S <= "000000001001" + P_HR_S406;
				when "01111100010" => P_HR_S <= "000000001001" + P_HR_S407;
				when "01111100101" => P_HR_S <= "000000010010" + P_HR_S408;
				when "01111101000" => P_HR_S <= "000000001001" + P_HR_S409;
				when "01111101011" => P_HR_S <= "000000011010" + P_HR_S410;
				when "01111101110" => P_HR_S <= "000000010010" + P_HR_S411;
				when "01111110111" => P_HR_S <= "000000011010" + P_HR_S412;
				when "01111111101" => P_HR_S <= "000000100011" + P_HR_S413;
				when "10000000000" => P_HR_S <= "000000001001" + P_HR_S414;
				when "10000000100" => P_HR_S <= "000000001001" + P_HR_S415;
				when "10000000111" => P_HR_S <= "000000010010" + P_HR_S416;
				when "10000001010" => P_HR_S <= "000000011010" + P_HR_S417;
				when "10000001101" => P_HR_S <= "000000001001" + P_HR_S418;
				when "10000010000" => P_HR_S <= "000000100011" + P_HR_S419;
				when "10000010011" => P_HR_S <= "000000011010" + P_HR_S420;
				when "10000010111" => P_HR_S <= "000000011010" + P_HR_S421;
				when "10000011010" => P_HR_S <= "000000100011" + P_HR_S422;
				when "10000011101" => P_HR_S <= "000000100011" + P_HR_S423;
				when "10000100100" => P_HR_S <= "000000010010" + P_HR_S424;
				when "10000101011" => P_HR_S <= "000000011010" + P_HR_S425;
				when "10000101110" => P_HR_S <= "000000010010" + P_HR_S426;
				when "10000110001" => P_HR_S <= "000000001001" + P_HR_S427;
				when "10000111000" => P_HR_S <= "000000001001" + P_HR_S428;
				when others        => P_HR_S <= "000000000001";
			end case;
			stress_score <= P_TEMP_S * P_STRESS * P_EDA_S * P_HR_S;
		
        -- score calc
		--stress_score <= P_TEMP_S * P_STRESS * P_EDA_S * P_HR_S;
		
		elsif state = TRAINING_S then
			
			case temp is
				when "011110111" =>P_TEMP_S1   <= P_TEMP_S1 + "01000";
				when "011111000" =>P_TEMP_S2   <= P_TEMP_S2 + "01000";
				when "011111001" =>P_TEMP_S3   <= P_TEMP_S3 + "01000";
				when "011111010" =>P_TEMP_S4   <= P_TEMP_S4 + "01000";
				when "011111011" =>P_TEMP_S5   <= P_TEMP_S5 + "01000";
				when "011111100" =>P_TEMP_S6   <= P_TEMP_S6 + "01000";
				when "011111101" =>P_TEMP_S7   <= P_TEMP_S7 + "01000";
				when "011111110" =>P_TEMP_S8   <= P_TEMP_S8 + "01000";
				when "011111111" =>P_TEMP_S9   <= P_TEMP_S9 + "01000";
				when "100000000" =>P_TEMP_S10 <= P_TEMP_S10 + "01000";
				when "100000001" =>P_TEMP_S11 <= P_TEMP_S11 + "01000";
				when "100000010" =>P_TEMP_S12 <= P_TEMP_S12 + "01000";
				when "100000011" =>P_TEMP_S13 <= P_TEMP_S13 + "01000";
				when "100000100" =>P_TEMP_S14 <= P_TEMP_S14 + "01000";
				when "100000101" =>P_TEMP_S15 <= P_TEMP_S15 + "01000";
				when "100000110" =>P_TEMP_S16 <= P_TEMP_S16 + "01000";
				when "100000111" =>P_TEMP_S17 <= P_TEMP_S17 + "01000";
				when "100001000" =>P_TEMP_S18 <= P_TEMP_S18 + "01000";
				when "100001001" =>P_TEMP_S19 <= P_TEMP_S19 + "01000";
				when "100001010" =>P_TEMP_S20 <= P_TEMP_S20 + "01000";
				when "100001011" =>P_TEMP_S21 <= P_TEMP_S21 + "01000";
				when "100001100" =>P_TEMP_S22 <= P_TEMP_S22 + "01000";
				when "100001101" =>P_TEMP_S23 <= P_TEMP_S23 + "01000";
				when "100001110" =>P_TEMP_S24 <= P_TEMP_S24 + "01000";
				when "100001111" =>P_TEMP_S25 <= P_TEMP_S25 + "01000";
				when "100010000" =>P_TEMP_S26 <= P_TEMP_S26 + "01000";
				when "100010001" =>P_TEMP_S27 <= P_TEMP_S27 + "01000";
				when "100010010" =>P_TEMP_S28 <= P_TEMP_S28 + "01000";
				when "100010011" =>P_TEMP_S29 <= P_TEMP_S29 + "01000";
				when "100010100" =>P_TEMP_S30 <= P_TEMP_S30 + "01000";
				when  others     => null;
				
			end case;	
		
			case hr is
				when "00000001100" => P_HR_S1     <= P_HR_S1 + "1000";
				when "00000001110" => P_HR_S2     <= P_HR_S2 + "1000";
				when "00000010011" => P_HR_S3     <= P_HR_S3 + "1000";
				when "00000010111" => P_HR_S4     <= P_HR_S4 + "1000";
				when "00000011001" => P_HR_S5     <= P_HR_S5 + "1000";
				when "00000011100" => P_HR_S6     <= P_HR_S6 + "1000";
				when "00000100101" => P_HR_S7     <= P_HR_S7 + "1000";
				when "00000100110" => P_HR_S8     <= P_HR_S8 + "1000";
				when "00000110001" => P_HR_S9     <= P_HR_S9 + "1000";
				when "00001000111" => P_HR_S10   <= P_HR_S10 + "1000";
				when "00001001100" => P_HR_S11   <= P_HR_S11 + "1000";
				when "00001001101" => P_HR_S12   <= P_HR_S12 + "1000";
				when "00001001110" => P_HR_S13   <= P_HR_S13 + "1000";
				when "00001010001" => P_HR_S14   <= P_HR_S14 + "1000";
				when "00001010101" => P_HR_S15   <= P_HR_S15 + "1000";
				when "00001010111" => P_HR_S16   <= P_HR_S16 + "1000";
				when "00001011001" => P_HR_S17   <= P_HR_S17 + "1000";
				when "00001100001" => P_HR_S18   <= P_HR_S18 + "1000";
				when "00001100010" => P_HR_S19   <= P_HR_S19 + "1000";
				when "00001100011" => P_HR_S20   <= P_HR_S20 + "1000";
				when "00001110000" => P_HR_S21   <= P_HR_S21 + "1000";
				when "00001110001" => P_HR_S22   <= P_HR_S22 + "1000";
				when "00001110101" => P_HR_S23   <= P_HR_S23 + "1000";
				when "00001111000" => P_HR_S24   <= P_HR_S24 + "1000";
				when "00001111100" => P_HR_S25   <= P_HR_S25 + "1000";
				when "00001111111" => P_HR_S26   <= P_HR_S26 + "1000";
				when "00010000011" => P_HR_S27   <= P_HR_S27 + "1000";
				when "00010000111" => P_HR_S28   <= P_HR_S28 + "1000";
				when "00010001011" => P_HR_S29   <= P_HR_S29 + "1000";
				when "00010001110" => P_HR_S30   <= P_HR_S30 + "1000";
				when "00010001111" => P_HR_S31   <= P_HR_S31 + "1000";
				when "00010010000" => P_HR_S32   <= P_HR_S32 + "1000";
				when "00010010010" => P_HR_S33   <= P_HR_S33 + "1000";
				when "00010010011" => P_HR_S34   <= P_HR_S34 + "1000";
				when "00010010100" => P_HR_S35   <= P_HR_S35 + "1000";
				when "00010010101" => P_HR_S36   <= P_HR_S36 + "1000";
				when "00010011000" => P_HR_S37   <= P_HR_S37 + "1000";
				when "00010011110" => P_HR_S38   <= P_HR_S38 + "1000";
				when "00010100010" => P_HR_S39   <= P_HR_S39 + "1000";
				when "00010110101" => P_HR_S40   <= P_HR_S40 + "1000";
				when "00010110110" => P_HR_S41   <= P_HR_S41 + "1000";
				when "00010111000" => P_HR_S42   <= P_HR_S42 + "1000";
				when "00010111001" => P_HR_S43   <= P_HR_S43 + "1000";
				when "00010111100" => P_HR_S44   <= P_HR_S44 + "1000";
				when "00010111101" => P_HR_S45   <= P_HR_S45 + "1000";
				when "00010111110" => P_HR_S46   <= P_HR_S46 + "1000";
				when "00010111111" => P_HR_S47   <= P_HR_S47 + "1000";
				when "00011000000" => P_HR_S48   <= P_HR_S48 + "1000";
				when "00011000001" => P_HR_S49   <= P_HR_S49 + "1000";
				when "00011000101" => P_HR_S50   <= P_HR_S50 + "1000";
				when "00011000110" => P_HR_S51   <= P_HR_S51 + "1000";
				when "00011000111" => P_HR_S52   <= P_HR_S52 + "1000";
				when "00011001000" => P_HR_S53   <= P_HR_S53 + "1000";
				when "00011001001" => P_HR_S54   <= P_HR_S54 + "1000";
				when "00011001010" => P_HR_S55   <= P_HR_S55 + "1000";
				when "00011001011" => P_HR_S56   <= P_HR_S56 + "1000";
				when "00011001101" => P_HR_S57   <= P_HR_S57 + "1000";
				when "00011001110" => P_HR_S58   <= P_HR_S58 + "1000";
				when "00011010000" => P_HR_S59   <= P_HR_S59 + "1000";
				when "00011010001" => P_HR_S60   <= P_HR_S60 + "1000";
				when "00011010100" => P_HR_S61   <= P_HR_S61 + "1000";
				when "00011011010" => P_HR_S62   <= P_HR_S62 + "1000";
				when "00011100100" => P_HR_S63   <= P_HR_S63 + "1000";
				when "00011111001" => P_HR_S64   <= P_HR_S64 + "1000";
				when "00100001111" => P_HR_S65   <= P_HR_S65 + "1000";
				when "00100010000" => P_HR_S66   <= P_HR_S66 + "1000";
				when "00100010001" => P_HR_S67   <= P_HR_S67 + "1000";
				when "00100010100" => P_HR_S68   <= P_HR_S68 + "1000";
				when "00100011001" => P_HR_S69   <= P_HR_S69 + "1000";
				when "00100011011" => P_HR_S70   <= P_HR_S70 + "1000";
				when "00100011100" => P_HR_S71   <= P_HR_S71 + "1000";
				when "00100011110" => P_HR_S72   <= P_HR_S72 + "1000";
				when "00100011111" => P_HR_S73   <= P_HR_S73 + "1000";
				when "00100100000" => P_HR_S74   <= P_HR_S74 + "1000";
				when "00100100001" => P_HR_S75   <= P_HR_S75 + "1000";
				when "00100100010" => P_HR_S76   <= P_HR_S76 + "1000";
				when "00100100011" => P_HR_S77   <= P_HR_S77 + "1000";
				when "00100100100" => P_HR_S78   <= P_HR_S78 + "1000";
				when "00100100101" => P_HR_S79   <= P_HR_S79 + "1000";
				when "00100100110" => P_HR_S80   <= P_HR_S80 + "1000";
				when "00100100111" => P_HR_S81   <= P_HR_S81 + "1000";
				when "00100101010" => P_HR_S82   <= P_HR_S82 + "1000";
				when "00100101100" => P_HR_S83   <= P_HR_S83 + "1000";
				when "00100101110" => P_HR_S84   <= P_HR_S84 + "1000";
				when "00100110010" => P_HR_S85   <= P_HR_S85 + "1000";
				when "00100110011" => P_HR_S86   <= P_HR_S86 + "1000";
				when "00100110100" => P_HR_S87   <= P_HR_S87 + "1000";
				when "00100110111" => P_HR_S88   <= P_HR_S88 + "1000";
				when "00100111000" => P_HR_S89   <= P_HR_S89 + "1000";
				when "00100111001" => P_HR_S90   <= P_HR_S90 + "1000";
				when "00100111101" => P_HR_S91   <= P_HR_S91 + "1000";
				when "00101000101" => P_HR_S92   <= P_HR_S92 + "1000";
				when "00101001101" => P_HR_S93   <= P_HR_S93 + "1000";
				when "00101010010" => P_HR_S94   <= P_HR_S94 + "1000";
				when "00101010100" => P_HR_S95   <= P_HR_S95 + "1000";
				when "00101011001" => P_HR_S96   <= P_HR_S96 + "1000";
				when "00110010011" => P_HR_S97   <= P_HR_S97 + "1000";
				when "00110010111" => P_HR_S98   <= P_HR_S98 + "1000";
				when "00110011000" => P_HR_S99   <= P_HR_S99 + "1000";
				when "00110011001" => P_HR_S100 <= P_HR_S100 + "1000";
				when "00110110011" => P_HR_S101 <= P_HR_S101 + "1000";
				when "00110110110" => P_HR_S102 <= P_HR_S102 + "1000";
				when "00110111100" => P_HR_S103 <= P_HR_S103 + "1000";
				when "00110111110" => P_HR_S104 <= P_HR_S104 + "1000";
				when "00111000000" => P_HR_S105 <= P_HR_S105 + "1000";
				when "00111000010" => P_HR_S106 <= P_HR_S106 + "1000";
				when "00111000011" => P_HR_S107 <= P_HR_S107 + "1000";
				when "00111000111" => P_HR_S108 <= P_HR_S108 + "1000";
				when "00111001001" => P_HR_S109 <= P_HR_S109 + "1000";
				when "00111001100" => P_HR_S110 <= P_HR_S110 + "1000";
				when "00111001101" => P_HR_S111 <= P_HR_S111 + "1000";
				when "00111001111" => P_HR_S112 <= P_HR_S112 + "1000";
				when "00111010010" => P_HR_S113 <= P_HR_S113 + "1000";
				when "00111010101" => P_HR_S114 <= P_HR_S114 + "1000";
				when "00111010111" => P_HR_S115 <= P_HR_S115 + "1000";
				when "00111011000" => P_HR_S116 <= P_HR_S116 + "1000";
				when "00111011001" => P_HR_S117 <= P_HR_S117 + "1000";
				when "00111011100" => P_HR_S118 <= P_HR_S118 + "1000";
				when "00111011101" => P_HR_S119 <= P_HR_S119 + "1000";
				when "00111100001" => P_HR_S120 <= P_HR_S120 + "1000";
				when "00111100011" => P_HR_S121 <= P_HR_S121 + "1000";
				when "00111100110" => P_HR_S122 <= P_HR_S122 + "1000";
				when "00111101011" => P_HR_S123 <= P_HR_S123 + "1000";
				when "00111101111" => P_HR_S124 <= P_HR_S124 + "1000";
				when "00111110000" => P_HR_S125 <= P_HR_S125 + "1000";
				when "00111110010" => P_HR_S126 <= P_HR_S126 + "1000";
				when "00111110100" => P_HR_S127 <= P_HR_S127 + "1000";
				when "00111110101" => P_HR_S128 <= P_HR_S128 + "1000";
				when "00111110110" => P_HR_S129 <= P_HR_S129 + "1000";
				when "00111111000" => P_HR_S130 <= P_HR_S130 + "1000";
				when "00111111001" => P_HR_S131 <= P_HR_S131 + "1000";
				when "00111111100" => P_HR_S132 <= P_HR_S132 + "1000";
				when "00111111111" => P_HR_S133 <= P_HR_S133 + "1000";
				when "01000000011" => P_HR_S134 <= P_HR_S134 + "1000";
				when "01000000100" => P_HR_S135 <= P_HR_S135 + "1000";
				when "01000000101" => P_HR_S136 <= P_HR_S136 + "1000";
				when "01000000110" => P_HR_S137 <= P_HR_S137 + "1000";
				when "01000000111" => P_HR_S138 <= P_HR_S138 + "1000";
				when "01000001001" => P_HR_S139 <= P_HR_S139 + "1000";
				when "01000001010" => P_HR_S140 <= P_HR_S140 + "1000";
				when "01000001011" => P_HR_S141 <= P_HR_S141 + "1000";
				when "01000001101" => P_HR_S142 <= P_HR_S142 + "1000";
				when "01000001111" => P_HR_S143 <= P_HR_S143 + "1000";
				when "01000010001" => P_HR_S144 <= P_HR_S144 + "1000";
				when "01000010010" => P_HR_S145 <= P_HR_S145 + "1000";
				when "01000010100" => P_HR_S146 <= P_HR_S146 + "1000";
				when "01000010101" => P_HR_S147 <= P_HR_S147 + "1000";
				when "01000010110" => P_HR_S148 <= P_HR_S148 + "1000";
				when "01000010111" => P_HR_S149 <= P_HR_S149 + "1000";
				when "01000011000" => P_HR_S150 <= P_HR_S150 + "1000";
				when "01000011010" => P_HR_S151 <= P_HR_S151 + "1000";
				when "01000011011" => P_HR_S152 <= P_HR_S152 + "1000";
				when "01000011100" => P_HR_S153 <= P_HR_S153 + "1000";
				when "01000011101" => P_HR_S154 <= P_HR_S154 + "1000";
				when "01000011111" => P_HR_S155 <= P_HR_S155 + "1000";
				when "01000100000" => P_HR_S156 <= P_HR_S156 + "1000";
				when "01000100001" => P_HR_S157 <= P_HR_S157 + "1000";
				when "01000100011" => P_HR_S158 <= P_HR_S158 + "1000";
				when "01000100100" => P_HR_S159 <= P_HR_S159 + "1000";
				when "01000100111" => P_HR_S160 <= P_HR_S160 + "1000";
				when "01000101000" => P_HR_S161 <= P_HR_S161 + "1000";
				when "01000101001" => P_HR_S162 <= P_HR_S162 + "1000";
				when "01000101010" => P_HR_S163 <= P_HR_S163 + "1000";
				when "01000101011" => P_HR_S164 <= P_HR_S164 + "1000";
				when "01000101100" => P_HR_S165 <= P_HR_S165 + "1000";
				when "01000101101" => P_HR_S166 <= P_HR_S166 + "1000";
				when "01000101110" => P_HR_S167 <= P_HR_S167 + "1000";
				when "01000101111" => P_HR_S168 <= P_HR_S168 + "1000";
				when "01000110000" => P_HR_S169 <= P_HR_S169 + "1000";
				when "01000110001" => P_HR_S170 <= P_HR_S170 + "1000";
				when "01000110011" => P_HR_S171 <= P_HR_S171 + "1000";
				when "01000110100" => P_HR_S172 <= P_HR_S172 + "1000";
				when "01000110101" => P_HR_S173 <= P_HR_S173 + "1000";
				when "01000110110" => P_HR_S174 <= P_HR_S174 + "1000";
				when "01000110111" => P_HR_S175 <= P_HR_S175 + "1000";
				when "01000111000" => P_HR_S176 <= P_HR_S176 + "1000";
				when "01000111001" => P_HR_S177 <= P_HR_S177 + "1000";
				when "01000111010" => P_HR_S178 <= P_HR_S178 + "1000";
				when "01000111011" => P_HR_S179 <= P_HR_S179 + "1000";
				when "01000111100" => P_HR_S180 <= P_HR_S180 + "1000";
				when "01000111101" => P_HR_S181 <= P_HR_S181 + "1000";
				when "01000111110" => P_HR_S182 <= P_HR_S182 + "1000";
				when "01000111111" => P_HR_S183 <= P_HR_S183 + "1000";
				when "01001000000" => P_HR_S184 <= P_HR_S184 + "1000";
				when "01001000001" => P_HR_S185 <= P_HR_S185 + "1000";
				when "01001000010" => P_HR_S186 <= P_HR_S186 + "1000";
				when "01001000011" => P_HR_S187 <= P_HR_S187 + "1000";
				when "01001000100" => P_HR_S188 <= P_HR_S188 + "1000";
				when "01001000101" => P_HR_S189 <= P_HR_S189 + "1000";
				when "01001000110" => P_HR_S190 <= P_HR_S190 + "1000";
				when "01001000111" => P_HR_S191 <= P_HR_S191 + "1000";
				when "01001001000" => P_HR_S192 <= P_HR_S192 + "1000";
				when "01001001001" => P_HR_S193 <= P_HR_S193 + "1000";
				when "01001001010" => P_HR_S194 <= P_HR_S194 + "1000";
				when "01001001011" => P_HR_S195 <= P_HR_S195 + "1000";
				when "01001001100" => P_HR_S196 <= P_HR_S196 + "1000";
				when "01001001101" => P_HR_S197 <= P_HR_S197 + "1000";
				when "01001001111" => P_HR_S198 <= P_HR_S198 + "1000";
				when "01001010001" => P_HR_S199 <= P_HR_S199 + "1000";
				when "01001010010" => P_HR_S200 <= P_HR_S200 + "1000";
				when "01001010011" => P_HR_S201 <= P_HR_S201 + "1000";
				when "01001010100" => P_HR_S202 <= P_HR_S202 + "1000";
				when "01001010101" => P_HR_S203 <= P_HR_S203 + "1000";
				when "01001010110" => P_HR_S204 <= P_HR_S204 + "1000";
				when "01001010111" => P_HR_S205 <= P_HR_S205 + "1000";
				when "01001011000" => P_HR_S206 <= P_HR_S206 + "1000";
				when "01001011001" => P_HR_S207 <= P_HR_S207 + "1000";
				when "01001011010" => P_HR_S208 <= P_HR_S208 + "1000";
				when "01001011011" => P_HR_S209 <= P_HR_S209 + "1000";
				when "01001011100" => P_HR_S210 <= P_HR_S210 + "1000";
				when "01001011101" => P_HR_S211 <= P_HR_S211 + "1000";
				when "01001011110" => P_HR_S212 <= P_HR_S212 + "1000";
				when "01001100001" => P_HR_S213 <= P_HR_S213 + "1000";
				when "01001100010" => P_HR_S214 <= P_HR_S214 + "1000";
				when "01001100011" => P_HR_S215 <= P_HR_S215 + "1000";
				when "01001100100" => P_HR_S216 <= P_HR_S216 + "1000";
				when "01001100101" => P_HR_S217 <= P_HR_S217 + "1000";
				when "01001100110" => P_HR_S218 <= P_HR_S218 + "1000";
				when "01001100111" => P_HR_S219 <= P_HR_S219 + "1000";
				when "01001101001" => P_HR_S220 <= P_HR_S220 + "1000";
				when "01001101010" => P_HR_S221 <= P_HR_S221 + "1000";
				when "01001101011" => P_HR_S222 <= P_HR_S222 + "1000";
				when "01001101100" => P_HR_S223 <= P_HR_S223 + "1000";
				when "01001101101" => P_HR_S224 <= P_HR_S224 + "1000";
				when "01001101110" => P_HR_S225 <= P_HR_S225 + "1000";
				when "01001101111" => P_HR_S226 <= P_HR_S226 + "1000";
				when "01001110001" => P_HR_S227 <= P_HR_S227 + "1000";
				when "01001110011" => P_HR_S228 <= P_HR_S228 + "1000";
				when "01001110100" => P_HR_S229 <= P_HR_S229 + "1000";
				when "01001110101" => P_HR_S230 <= P_HR_S230 + "1000";
				when "01001110110" => P_HR_S231 <= P_HR_S231 + "1000";
				when "01001111000" => P_HR_S232 <= P_HR_S232 + "1000";
				when "01001111001" => P_HR_S233 <= P_HR_S233 + "1000";
				when "01001111010" => P_HR_S234 <= P_HR_S234 + "1000";
				when "01001111011" => P_HR_S235 <= P_HR_S235 + "1000";
				when "01001111100" => P_HR_S236 <= P_HR_S236 + "1000";
				when "01001111110" => P_HR_S237 <= P_HR_S237 + "1000";
				when "01001111111" => P_HR_S238 <= P_HR_S238 + "1000";
				when "01010000000" => P_HR_S239 <= P_HR_S239 + "1000";
				when "01010000001" => P_HR_S240 <= P_HR_S240 + "1000";
				when "01010000010" => P_HR_S241 <= P_HR_S241 + "1000";
				when "01010000100" => P_HR_S242 <= P_HR_S242 + "1000";
				when "01010000101" => P_HR_S243 <= P_HR_S243 + "1000";
				when "01010000110" => P_HR_S244 <= P_HR_S244 + "1000";
				when "01010001001" => P_HR_S245 <= P_HR_S245 + "1000";
				when "01010001010" => P_HR_S246 <= P_HR_S246 + "1000";
				when "01010001011" => P_HR_S247 <= P_HR_S247 + "1000";
				when "01010001110" => P_HR_S248 <= P_HR_S248 + "1000";
				when "01010001111" => P_HR_S249 <= P_HR_S249 + "1000";
				when "01010010000" => P_HR_S250 <= P_HR_S250 + "1000";
				when "01010010010" => P_HR_S251 <= P_HR_S251 + "1000";
				when "01010010011" => P_HR_S252 <= P_HR_S252 + "1000";
				when "01010010100" => P_HR_S253 <= P_HR_S253 + "1000";
				when "01010010101" => P_HR_S254 <= P_HR_S254 + "1000";
				when "01010010111" => P_HR_S255 <= P_HR_S255 + "1000";
				when "01010011000" => P_HR_S256 <= P_HR_S256 + "1000";
				when "01010011001" => P_HR_S257 <= P_HR_S257 + "1000";
				when "01010011011" => P_HR_S258 <= P_HR_S258 + "1000";
				when "01010011100" => P_HR_S259 <= P_HR_S259 + "1000";
				when "01010011101" => P_HR_S260 <= P_HR_S260 + "1000";
				when "01010011111" => P_HR_S261 <= P_HR_S261 + "1000";
				when "01010100000" => P_HR_S262 <= P_HR_S262 + "1000";
				when "01010100001" => P_HR_S263 <= P_HR_S263 + "1000";
				when "01010100011" => P_HR_S264 <= P_HR_S264 + "1000";
				when "01010100100" => P_HR_S265 <= P_HR_S265 + "1000";
				when "01010100101" => P_HR_S266 <= P_HR_S266 + "1000";
				when "01010100111" => P_HR_S267 <= P_HR_S267 + "1000";
				when "01010101000" => P_HR_S268 <= P_HR_S268 + "1000";
				when "01010101010" => P_HR_S269 <= P_HR_S269 + "1000";
				when "01010101011" => P_HR_S270 <= P_HR_S270 + "1000";
				when "01010101100" => P_HR_S271 <= P_HR_S271 + "1000";
				when "01010101110" => P_HR_S272 <= P_HR_S272 + "1000";
				when "01010101111" => P_HR_S273 <= P_HR_S273 + "1000";
				when "01010110001" => P_HR_S274 <= P_HR_S274 + "1000";
				when "01010110010" => P_HR_S275 <= P_HR_S275 + "1000";
				when "01010110011" => P_HR_S276 <= P_HR_S276 + "1000";
				when "01010110101" => P_HR_S277 <= P_HR_S277 + "1000";
				when "01010110110" => P_HR_S278 <= P_HR_S278 + "1000";
				when "01010111000" => P_HR_S279 <= P_HR_S279 + "1000";
				when "01010111001" => P_HR_S280 <= P_HR_S280 + "1000";
				when "01010111100" => P_HR_S281 <= P_HR_S281 + "1000";
				when "01010111101" => P_HR_S282 <= P_HR_S282 + "1000";
				when "01010111111" => P_HR_S283 <= P_HR_S283 + "1000";
				when "01011000000" => P_HR_S284 <= P_HR_S284 + "1000";
				when "01011000010" => P_HR_S285 <= P_HR_S285 + "1000";
				when "01011000011" => P_HR_S286 <= P_HR_S286 + "1000";
				when "01011000101" => P_HR_S287 <= P_HR_S287 + "1000";
				when "01011000110" => P_HR_S288 <= P_HR_S288 + "1000";
				when "01011001000" => P_HR_S289 <= P_HR_S289 + "1000";
				when "01011001001" => P_HR_S290 <= P_HR_S290 + "1000";
				when "01011001011" => P_HR_S291 <= P_HR_S291 + "1000";
				when "01011001100" => P_HR_S292 <= P_HR_S292 + "1000";
				when "01011001110" => P_HR_S293 <= P_HR_S293 + "1000";
				when "01011001111" => P_HR_S294 <= P_HR_S294 + "1000";
				when "01011010001" => P_HR_S295 <= P_HR_S295 + "1000";
				when "01011010011" => P_HR_S296 <= P_HR_S296 + "1000";
				when "01011010100" => P_HR_S297 <= P_HR_S297 + "1000";
				when "01011010110" => P_HR_S298 <= P_HR_S298 + "1000";
				when "01011010111" => P_HR_S299 <= P_HR_S299 + "1000";
				when "01011011001" => P_HR_S300 <= P_HR_S300 + "1000";
				when "01011011010" => P_HR_S301 <= P_HR_S301 + "1000";
				when "01011011100" => P_HR_S302 <= P_HR_S302 + "1000";
				when "01011011110" => P_HR_S303 <= P_HR_S303 + "1000";
				when "01011011111" => P_HR_S304 <= P_HR_S304 + "1000";
				when "01011100001" => P_HR_S305 <= P_HR_S305 + "1000";
				when "01011100010" => P_HR_S306 <= P_HR_S306 + "1000";
				when "01011100100" => P_HR_S307 <= P_HR_S307 + "1000";
				when "01011100110" => P_HR_S308 <= P_HR_S308 + "1000";
				when "01011100111" => P_HR_S309 <= P_HR_S309 + "1000";
				when "01011101001" => P_HR_S310 <= P_HR_S310 + "1000";
				when "01011101011" => P_HR_S311 <= P_HR_S311 + "1000";
				when "01011101100" => P_HR_S312 <= P_HR_S312 + "1000";
				when "01011101110" => P_HR_S313 <= P_HR_S313 + "1000";
				when "01011110000" => P_HR_S314 <= P_HR_S314 + "1000";
				when "01011110001" => P_HR_S315 <= P_HR_S315 + "1000";
				when "01011110011" => P_HR_S316 <= P_HR_S316 + "1000";
				when "01011110101" => P_HR_S317 <= P_HR_S317 + "1000";
				when "01011110110" => P_HR_S318 <= P_HR_S318 + "1000";
				when "01011111000" => P_HR_S319 <= P_HR_S319 + "1000";
				when "01011111010" => P_HR_S320 <= P_HR_S320 + "1000";
				when "01011111100" => P_HR_S321 <= P_HR_S321 + "1000";
				when "01011111101" => P_HR_S322 <= P_HR_S322 + "1000";
				when "01011111111" => P_HR_S323 <= P_HR_S323 + "1000";
				when "01100000001" => P_HR_S324 <= P_HR_S324 + "1000";
				when "01100000011" => P_HR_S325 <= P_HR_S325 + "1000";
				when "01100000100" => P_HR_S326 <= P_HR_S326 + "1000";
				when "01100000110" => P_HR_S327 <= P_HR_S327 + "1000";
				when "01100001000" => P_HR_S328 <= P_HR_S328 + "1000";
				when "01100001010" => P_HR_S329 <= P_HR_S329 + "1000";
				when "01100001100" => P_HR_S330 <= P_HR_S330 + "1000";
				when "01100001101" => P_HR_S331 <= P_HR_S331 + "1000";
				when "01100001111" => P_HR_S332 <= P_HR_S332 + "1000";
				when "01100010001" => P_HR_S333 <= P_HR_S333 + "1000";
				when "01100010011" => P_HR_S334 <= P_HR_S334 + "1000";
				when "01100010101" => P_HR_S335 <= P_HR_S335 + "1000";
				when "01100010111" => P_HR_S336 <= P_HR_S336 + "1000";
				when "01100011000" => P_HR_S337 <= P_HR_S337 + "1000";
				when "01100011010" => P_HR_S338 <= P_HR_S338 + "1000";
				when "01100011110" => P_HR_S339 <= P_HR_S339 + "1000";
				when "01100100000" => P_HR_S340 <= P_HR_S340 + "1000";
				when "01100100010" => P_HR_S341 <= P_HR_S341 + "1000";
				when "01100100100" => P_HR_S342 <= P_HR_S342 + "1000";
				when "01100100110" => P_HR_S343 <= P_HR_S343 + "1000";
				when "01100101000" => P_HR_S344 <= P_HR_S344 + "1000";
				when "01100101010" => P_HR_S345 <= P_HR_S345 + "1000";
				when "01100101100" => P_HR_S346 <= P_HR_S346 + "1000";
				when "01100101110" => P_HR_S347 <= P_HR_S347 + "1000";
				when "01100110000" => P_HR_S348 <= P_HR_S348 + "1000";
				when "01100110010" => P_HR_S349 <= P_HR_S349 + "1000";
				when "01100110100" => P_HR_S350 <= P_HR_S350 + "1000";
				when "01100110110" => P_HR_S351 <= P_HR_S351 + "1000";
				when "01100111000" => P_HR_S352 <= P_HR_S352 + "1000";
				when "01100111010" => P_HR_S353 <= P_HR_S353 + "1000";
				when "01100111100" => P_HR_S354 <= P_HR_S354 + "1000";
				when "01100111110" => P_HR_S355 <= P_HR_S355 + "1000";
				when "01101000000" => P_HR_S356 <= P_HR_S356 + "1000";
				when "01101000010" => P_HR_S357 <= P_HR_S357 + "1000";
				when "01101000100" => P_HR_S358 <= P_HR_S358 + "1000";
				when "01101000110" => P_HR_S359 <= P_HR_S359 + "1000";
				when "01101001000" => P_HR_S360 <= P_HR_S360 + "1000";
				when "01101001100" => P_HR_S361 <= P_HR_S361 + "1000";
				when "01101001110" => P_HR_S362 <= P_HR_S362 + "1000";
				when "01101010000" => P_HR_S363 <= P_HR_S363 + "1000";
				when "01101010011" => P_HR_S364 <= P_HR_S364 + "1000";
				when "01101010101" => P_HR_S365 <= P_HR_S365 + "1000";
				when "01101010111" => P_HR_S366 <= P_HR_S366 + "1000";
				when "01101011001" => P_HR_S367 <= P_HR_S367 + "1000";
				when "01101011011" => P_HR_S368 <= P_HR_S368 + "1000";
				when "01101011110" => P_HR_S369 <= P_HR_S369 + "1000";
				when "01101100000" => P_HR_S370 <= P_HR_S370 + "1000";
				when "01101100010" => P_HR_S371 <= P_HR_S371 + "1000";
				when "01101100100" => P_HR_S372 <= P_HR_S372 + "1000";
				when "01101100110" => P_HR_S373 <= P_HR_S373 + "1000";
				when "01101101001" => P_HR_S374 <= P_HR_S374 + "1000";
				when "01101101011" => P_HR_S375 <= P_HR_S375 + "1000";
				when "01101101101" => P_HR_S376 <= P_HR_S376 + "1000";
				when "01101110000" => P_HR_S377 <= P_HR_S377 + "1000";
				when "01101110010" => P_HR_S378 <= P_HR_S378 + "1000";
				when "01101110100" => P_HR_S379 <= P_HR_S379 + "1000";
				when "01101111011" => P_HR_S380 <= P_HR_S380 + "1000";
				when "01101111110" => P_HR_S381 <= P_HR_S381 + "1000";
				when "01110000101" => P_HR_S382 <= P_HR_S382 + "1000";
				when "01110000111" => P_HR_S383 <= P_HR_S383 + "1000";
				when "01110001010" => P_HR_S384 <= P_HR_S384 + "1000";
				when "01110001100" => P_HR_S385 <= P_HR_S385 + "1000";
				when "01110001111" => P_HR_S386 <= P_HR_S386 + "1000";
				when "01110010100" => P_HR_S387 <= P_HR_S387 + "1000";
				when "01110010110" => P_HR_S388 <= P_HR_S388 + "1000";
				when "01110011001" => P_HR_S389 <= P_HR_S389 + "1000";
				when "01110011011" => P_HR_S390 <= P_HR_S390 + "1000";
				when "01110100011" => P_HR_S391 <= P_HR_S391 + "1000";
				when "01110101101" => P_HR_S392 <= P_HR_S392 + "1000";
				when "01110110010" => P_HR_S393 <= P_HR_S393 + "1000";
				when "01110110101" => P_HR_S394 <= P_HR_S394 + "1000";
				when "01110111000" => P_HR_S395 <= P_HR_S395 + "1000";
				when "01110111011" => P_HR_S396 <= P_HR_S396 + "1000";
				when "01111000000" => P_HR_S397 <= P_HR_S397 + "1000";
				when "01111000110" => P_HR_S398 <= P_HR_S398 + "1000";
				when "01111001000" => P_HR_S399 <= P_HR_S399 + "1000";
				when "01111001011" => P_HR_S400 <= P_HR_S400 + "1000";
				when "01111001110" => P_HR_S401 <= P_HR_S401 + "1000";
				when "01111010001" => P_HR_S402 <= P_HR_S402 + "1000";
				when "01111010100" => P_HR_S403 <= P_HR_S403 + "1000";
				when "01111010110" => P_HR_S404 <= P_HR_S404 + "1000";
				when "01111011100" => P_HR_S405 <= P_HR_S405 + "1000";
				when "01111011111" => P_HR_S406 <= P_HR_S406 + "1000";
				when "01111100010" => P_HR_S407 <= P_HR_S407 + "1000";
				when "01111100101" => P_HR_S408 <= P_HR_S408 + "1000";
				when "01111101000" => P_HR_S409 <= P_HR_S409 + "1000";
				when "01111101011" => P_HR_S410 <= P_HR_S410 + "1000";
				when "01111101110" => P_HR_S411 <= P_HR_S411 + "1000";
				when "01111110111" => P_HR_S412 <= P_HR_S412 + "1000";
				when "01111111101" => P_HR_S413 <= P_HR_S413 + "1000";
				when "10000000000" => P_HR_S414 <= P_HR_S414 + "1000";
				when "10000000100" => P_HR_S415 <= P_HR_S415 + "1000";
				when "10000000111" => P_HR_S416 <= P_HR_S416 + "1000";
				when "10000001010" => P_HR_S417 <= P_HR_S417 + "1000";
				when "10000001101" => P_HR_S418 <= P_HR_S418 + "1000";
				when "10000010000" => P_HR_S419 <= P_HR_S419 + "1000";
				when "10000010011" => P_HR_S420 <= P_HR_S420 + "1000";
				when "10000010111" => P_HR_S421 <= P_HR_S421 + "1000";
				when "10000011010" => P_HR_S422 <= P_HR_S422 + "1000";
				when "10000011101" => P_HR_S423 <= P_HR_S423 + "1000";
				when "10000100100" => P_HR_S424 <= P_HR_S424 + "1000";
				when "10000101011" => P_HR_S425 <= P_HR_S425 + "1000";
				when "10000101110" => P_HR_S426 <= P_HR_S426 + "1000";
				when "10000110001" => P_HR_S427 <= P_HR_S427 + "1000";
				when "10000111000" => P_HR_S428 <= P_HR_S428 + "1000";
				when others            => null;
			end case;

			case eda is
			    when "0001000" => P_EDA_S1   <= P_EDA_S1 + "1000";
				when "0001001" => P_EDA_S2   <= P_EDA_S2 + "1000";
				when "0001010" => P_EDA_S3   <= P_EDA_S3 + "1000";
				when "0001011" => P_EDA_S4   <= P_EDA_S4 + "1000";
				when "0001100" => P_EDA_S5   <= P_EDA_S5 + "1000";
				when "0001101" => P_EDA_S6   <= P_EDA_S6 + "1000";
				when "0001110" => P_EDA_S7   <= P_EDA_S7 + "1000";
				when "0001111" => P_EDA_S8   <= P_EDA_S8 + "1000";
				when "0010000" => P_EDA_S9   <= P_EDA_S9 + "1000";
				when "0010001" => P_EDA_S10 <= P_EDA_S10 + "1000";
				when "0010010" => P_EDA_S11 <= P_EDA_S11 + "1000";
				when "0010011" => P_EDA_S12 <= P_EDA_S12 + "1000";
				when "0010100" => P_EDA_S13 <= P_EDA_S13 + "1000";
				when "0010101" => P_EDA_S14 <= P_EDA_S14 + "1000";
				when "0010110" => P_EDA_S15 <= P_EDA_S15 + "1000";
				when "0010111" => P_EDA_S16 <= P_EDA_S16 + "1000";
				when "0011000" => P_EDA_S17 <= P_EDA_S17 + "1000";
				when "0011001" => P_EDA_S18 <= P_EDA_S18 + "1000";
				when "0011010" => P_EDA_S19 <= P_EDA_S19 + "1000";
				when "0011011" => P_EDA_S20 <= P_EDA_S20 + "1000";
				when "0011100" => P_EDA_S21 <= P_EDA_S21 + "1000";
				when "0110110" => P_EDA_S22 <= P_EDA_S22 + "1000";
				when "0110111" => P_EDA_S23 <= P_EDA_S23 + "1000";
				when "0111000" => P_EDA_S24 <= P_EDA_S24 + "1000";
				when "0111001" => P_EDA_S25 <= P_EDA_S25 + "1000";
				when "0111010" => P_EDA_S26 <= P_EDA_S26 + "1000";
				when "0111011" => P_EDA_S27 <= P_EDA_S27 + "1000";
				when "0111100" => P_EDA_S28 <= P_EDA_S28 + "1000";
				when "0111101" => P_EDA_S29 <= P_EDA_S29 + "1000";
				when "0111110" => P_EDA_S30 <= P_EDA_S30 + "1000";
				when "0111111" => P_EDA_S31 <= P_EDA_S31 + "1000";
				when "1000000" => P_EDA_S32 <= P_EDA_S32 + "1000";
				when "1000001" => P_EDA_S33 <= P_EDA_S33 + "1000";
				when "1000010" => P_EDA_S34 <= P_EDA_S34 + "1000";
				when "1000011" => P_EDA_S35 <= P_EDA_S35 + "1000";
				when "1000100" => P_EDA_S36 <= P_EDA_S36 + "1000";
				when "1000101" => P_EDA_S37 <= P_EDA_S37 + "1000";
				when "1000110" => P_EDA_S38 <= P_EDA_S38 + "1000";
				when "1000111" => P_EDA_S39 <= P_EDA_S39 + "1000";
				when "1001000" => P_EDA_S40 <= P_EDA_S40 + "1000";
				when "1001001" => P_EDA_S41 <= P_EDA_S41 + "1000";
				when "1001010" => P_EDA_S42 <= P_EDA_S42 + "1000";
				when "1001011" => P_EDA_S43 <= P_EDA_S43 + "1000";
				when "1001100" => P_EDA_S44 <= P_EDA_S44 + "1000";
				when "1001101" => P_EDA_S45 <= P_EDA_S45 + "1000";
				when "1001110" => P_EDA_S46 <= P_EDA_S46 + "1000";
				when "1001111" => P_EDA_S47 <= P_EDA_S47 + "1000";
				when "1010000" => P_EDA_S48 <= P_EDA_S48 + "1000";
				when "1010001" => P_EDA_S49 <= P_EDA_S49 + "1000";
				when "1010010" => P_EDA_S50 <= P_EDA_S50 + "1000";
				when "1010011" => P_EDA_S51 <= P_EDA_S51 + "1000";
				when "1010100" => P_EDA_S52 <= P_EDA_S52 + "1000";
				when "1010101" => P_EDA_S53 <= P_EDA_S53 + "1000";
				when "1010110" => P_EDA_S54 <= P_EDA_S54 + "1000";
				when "1010111" => P_EDA_S55 <= P_EDA_S55 + "1000";
				when "1011000" => P_EDA_S56 <= P_EDA_S56 + "1000";
				when "1011001" => P_EDA_S57 <= P_EDA_S57 + "1000";
				when "1011010" => P_EDA_S58 <= P_EDA_S58 + "1000";
				when "1011011" => P_EDA_S59 <= P_EDA_S59 + "1000";
				when "1011100" => P_EDA_S60 <= P_EDA_S60 + "1000";
				when "1011101" => P_EDA_S61 <= P_EDA_S61 + "1000";
				when "1011110" => P_EDA_S62 <= P_EDA_S62 + "1000";
				when "1011111" => P_EDA_S63 <= P_EDA_S63 + "1000";
				when "1100000" => P_EDA_S64 <= P_EDA_S64 + "1000";
				when "1100001" => P_EDA_S65 <= P_EDA_S65 + "1000";
				when others            => null;
			end case;
		    
		else -- in training mode
			stress_score <= (others => '0');
			P_TEMP_S <= (others => '0'); 
			P_EDA_S <= (others => '0');
			P_HR_S <= (others => '0');
		end if;
		end if;
	end process;
	
	process(clk, rst) -- not stressed
	begin
	if (rst = '1') then
		-- reset logic
		P_TEMP_NS1 <= (others => '0');
		P_TEMP_NS2 <= (others => '0');
		P_TEMP_NS3 <= (others => '0');
		P_TEMP_NS4 <= (others => '0');
		P_TEMP_NS5 <= (others => '0');
		P_TEMP_NS6 <= (others => '0');
		P_TEMP_NS7 <= (others => '0');
		P_TEMP_NS8 <= (others => '0');
		P_TEMP_NS9 <= (others => '0');
		P_TEMP_NS10 <= (others => '0');
		P_TEMP_NS11 <= (others => '0');
		P_TEMP_NS12 <= (others => '0');
		P_TEMP_NS13 <= (others => '0');
		P_TEMP_NS14 <= (others => '0');
		P_TEMP_NS15 <= (others => '0');
		P_TEMP_NS16 <= (others => '0');
		P_TEMP_NS17 <= (others => '0');
		P_TEMP_NS18 <= (others => '0');
		P_TEMP_NS19 <= (others => '0');
		P_TEMP_NS20 <= (others => '0');
		P_TEMP_NS21 <= (others => '0');
		P_TEMP_NS22 <= (others => '0');
		P_TEMP_NS23 <= (others => '0');
		P_TEMP_NS24 <= (others => '0');
		P_TEMP_NS25 <= (others => '0');
		P_TEMP_NS26 <= (others => '0');
		P_TEMP_NS27 <= (others => '0');
		P_TEMP_NS28 <= (others => '0');
		P_TEMP_NS29 <= (others => '0');
		P_TEMP_NS30 <= (others => '0');
		P_TEMP_NS31 <= (others => '0');
		P_TEMP_NS32 <= (others => '0');
		P_TEMP_NS33 <= (others => '0');
		P_TEMP_NS34 <= (others => '0');
		P_TEMP_NS35 <= (others => '0');
		P_TEMP_NS36 <= (others => '0');
		P_TEMP_NS37 <= (others => '0');
		P_TEMP_NS38 <= (others => '0');
		P_TEMP_NS39 <= (others => '0');
		P_TEMP_NS40 <= (others => '0');
		P_TEMP_NS41 <= (others => '0');
		P_TEMP_NS42 <= (others => '0');
		P_TEMP_NS43 <= (others => '0');
		P_TEMP_NS44 <= (others => '0');
		P_TEMP_NS45 <= (others => '0');
		P_TEMP_NS46 <= (others => '0');
		P_TEMP_NS47 <= (others => '0');
		P_TEMP_NS48 <= (others => '0');
		P_TEMP_NS49 <= (others => '0');
		P_TEMP_NS50 <= (others => '0');
		P_TEMP_NS51 <= (others => '0');
		P_TEMP_NS52 <= (others => '0');	
			
		P_HR_NS1 <= (others => '0');
		P_HR_NS2 <= (others => '0');
		P_HR_NS3 <= (others => '0');
		P_HR_NS4 <= (others => '0');
		P_HR_NS5 <= (others => '0');
		P_HR_NS6 <= (others => '0');
		P_HR_NS7 <= (others => '0');
		P_HR_NS8 <= (others => '0');
		P_HR_NS9 <= (others => '0');
		P_HR_NS10 <= (others => '0');
		P_HR_NS11 <= (others => '0');
		P_HR_NS12 <= (others => '0');
		P_HR_NS13 <= (others => '0');
		P_HR_NS14 <= (others => '0');
		P_HR_NS15 <= (others => '0');
		P_HR_NS16 <= (others => '0');
		P_HR_NS17 <= (others => '0');
		P_HR_NS18 <= (others => '0');
		P_HR_NS19 <= (others => '0');
		P_HR_NS20 <= (others => '0');
		P_HR_NS21 <= (others => '0');
		P_HR_NS22 <= (others => '0');
		P_HR_NS23 <= (others => '0');
		P_HR_NS24 <= (others => '0');
		P_HR_NS25 <= (others => '0');
		P_HR_NS26 <= (others => '0');
		P_HR_NS27 <= (others => '0');
		P_HR_NS28 <= (others => '0');
		P_HR_NS29 <= (others => '0');
		P_HR_NS30 <= (others => '0');
		P_HR_NS31 <= (others => '0');
		P_HR_NS32 <= (others => '0');
		P_HR_NS33 <= (others => '0');
		P_HR_NS34 <= (others => '0');
		P_HR_NS35 <= (others => '0');
		P_HR_NS36 <= (others => '0');
		P_HR_NS37 <= (others => '0');
		P_HR_NS38 <= (others => '0');
		P_HR_NS39 <= (others => '0');
		P_HR_NS40 <= (others => '0');
		P_HR_NS41 <= (others => '0');
		P_HR_NS42 <= (others => '0');
		P_HR_NS43 <= (others => '0');
		P_HR_NS44 <= (others => '0');
		P_HR_NS45 <= (others => '0');
		P_HR_NS46 <= (others => '0');
		P_HR_NS47 <= (others => '0');
		P_HR_NS48 <= (others => '0');
		P_HR_NS49 <= (others => '0');
		P_HR_NS50 <= (others => '0');
		P_HR_NS51 <= (others => '0');
		P_HR_NS52 <= (others => '0');
		P_HR_NS53 <= (others => '0');
		P_HR_NS54 <= (others => '0');
		P_HR_NS55 <= (others => '0');
		P_HR_NS56 <= (others => '0');
		P_HR_NS57 <= (others => '0');
		P_HR_NS58 <= (others => '0');
		P_HR_NS59 <= (others => '0');
		P_HR_NS60 <= (others => '0');
		P_HR_NS61 <= (others => '0');
		P_HR_NS62 <= (others => '0');
		P_HR_NS63 <= (others => '0');
		P_HR_NS64 <= (others => '0');
		P_HR_NS65 <= (others => '0');
		P_HR_NS66 <= (others => '0');
		P_HR_NS67 <= (others => '0');
		P_HR_NS68 <= (others => '0');
		P_HR_NS69 <= (others => '0');
		P_HR_NS70 <= (others => '0');
		P_HR_NS71 <= (others => '0');
		P_HR_NS72 <= (others => '0');
		P_HR_NS73 <= (others => '0');
		P_HR_NS74 <= (others => '0');
		P_HR_NS75 <= (others => '0');
		P_HR_NS76 <= (others => '0');
		P_HR_NS77 <= (others => '0');
		P_HR_NS78 <= (others => '0');
		P_HR_NS79 <= (others => '0');
		P_HR_NS80 <= (others => '0');
		P_HR_NS81 <= (others => '0');
		P_HR_NS82 <= (others => '0');
		P_HR_NS83 <= (others => '0');
		P_HR_NS84 <= (others => '0');
		P_HR_NS85 <= (others => '0');
		P_HR_NS86 <= (others => '0');
		P_HR_NS87 <= (others => '0');
		P_HR_NS88 <= (others => '0');
		P_HR_NS89 <= (others => '0');
		P_HR_NS90 <= (others => '0');
		P_HR_NS91 <= (others => '0');
		P_HR_NS92 <= (others => '0');
		P_HR_NS93 <= (others => '0');
		P_HR_NS94 <= (others => '0');
		P_HR_NS95 <= (others => '0');
		P_HR_NS96 <= (others => '0');
		P_HR_NS97 <= (others => '0');
		P_HR_NS98 <= (others => '0');
		P_HR_NS99 <= (others => '0');
		P_HR_NS100 <= (others => '0');
		P_HR_NS101 <= (others => '0');
		P_HR_NS102 <= (others => '0');
		P_HR_NS103 <= (others => '0');
		P_HR_NS104 <= (others => '0');
		P_HR_NS105 <= (others => '0');
		P_HR_NS106 <= (others => '0');
		P_HR_NS107 <= (others => '0');
		P_HR_NS108 <= (others => '0');
		P_HR_NS109 <= (others => '0');
		P_HR_NS110 <= (others => '0');
		P_HR_NS111 <= (others => '0');
		P_HR_NS112 <= (others => '0');
		P_HR_NS113 <= (others => '0');
		P_HR_NS114 <= (others => '0');
		P_HR_NS115 <= (others => '0');
		P_HR_NS116 <= (others => '0');
		P_HR_NS117 <= (others => '0');
		P_HR_NS118 <= (others => '0');
		P_HR_NS119 <= (others => '0');
		P_HR_NS120 <= (others => '0');
		P_HR_NS121 <= (others => '0');
		P_HR_NS122 <= (others => '0');
		P_HR_NS123 <= (others => '0');
		P_HR_NS124 <= (others => '0');
		P_HR_NS125 <= (others => '0');
		P_HR_NS126 <= (others => '0');
		P_HR_NS127 <= (others => '0');
		P_HR_NS128 <= (others => '0');
		P_HR_NS129 <= (others => '0');
		P_HR_NS130 <= (others => '0');
		P_HR_NS131 <= (others => '0');
		P_HR_NS132 <= (others => '0');
		P_HR_NS133 <= (others => '0');
		P_HR_NS134 <= (others => '0');
		P_HR_NS135 <= (others => '0');
		P_HR_NS136 <= (others => '0');
		P_HR_NS137 <= (others => '0');
		P_HR_NS138 <= (others => '0');
		P_HR_NS139 <= (others => '0');
		P_HR_NS140 <= (others => '0');
		P_HR_NS141 <= (others => '0');
		P_HR_NS142 <= (others => '0');
		P_HR_NS143 <= (others => '0');
		P_HR_NS144 <= (others => '0');
		P_HR_NS145 <= (others => '0');
		P_HR_NS146 <= (others => '0');
		P_HR_NS147 <= (others => '0');
		P_HR_NS148 <= (others => '0');
		P_HR_NS149 <= (others => '0');
		P_HR_NS150 <= (others => '0');
		P_HR_NS151 <= (others => '0');
		P_HR_NS152 <= (others => '0');
		P_HR_NS153 <= (others => '0');
		P_HR_NS154 <= (others => '0');
		P_HR_NS155 <= (others => '0');
		P_HR_NS156 <= (others => '0');
		P_HR_NS157 <= (others => '0');
		P_HR_NS158 <= (others => '0');
		P_HR_NS159 <= (others => '0');
		P_HR_NS160 <= (others => '0');
		P_HR_NS161 <= (others => '0');
		P_HR_NS162 <= (others => '0');
		P_HR_NS163 <= (others => '0');
		P_HR_NS164 <= (others => '0');
		P_HR_NS165 <= (others => '0');
		P_HR_NS166 <= (others => '0');
		P_HR_NS167 <= (others => '0');
		P_HR_NS168 <= (others => '0');
		P_HR_NS169 <= (others => '0');
		P_HR_NS170 <= (others => '0');
		P_HR_NS171 <= (others => '0');
		P_HR_NS172 <= (others => '0');
		P_HR_NS173 <= (others => '0');
		P_HR_NS174 <= (others => '0');
		P_HR_NS175 <= (others => '0');
		P_HR_NS176 <= (others => '0');
		P_HR_NS177 <= (others => '0');
		P_HR_NS178 <= (others => '0');
		P_HR_NS179 <= (others => '0');
		P_HR_NS180 <= (others => '0');
		P_HR_NS181 <= (others => '0');
		P_HR_NS182 <= (others => '0');
		P_HR_NS183 <= (others => '0');
		P_HR_NS184 <= (others => '0');
		P_HR_NS185 <= (others => '0');
		P_HR_NS186 <= (others => '0');
		P_HR_NS187 <= (others => '0');
		P_HR_NS188 <= (others => '0');
		P_HR_NS189 <= (others => '0');
		P_HR_NS190 <= (others => '0');
		P_HR_NS191 <= (others => '0');
		P_HR_NS192 <= (others => '0');
		P_HR_NS193 <= (others => '0');
		P_HR_NS194 <= (others => '0');
		P_HR_NS195 <= (others => '0');
		P_HR_NS196 <= (others => '0');
		P_HR_NS197 <= (others => '0');
		P_HR_NS198 <= (others => '0');
		P_HR_NS199 <= (others => '0');
		P_HR_NS200 <= (others => '0');
		P_HR_NS201 <= (others => '0');
		P_HR_NS202 <= (others => '0');
		P_HR_NS203 <= (others => '0');
		P_HR_NS204 <= (others => '0');
		P_HR_NS205 <= (others => '0');
		P_HR_NS206 <= (others => '0');
		P_HR_NS207 <= (others => '0');
		P_HR_NS208 <= (others => '0');
		P_HR_NS209 <= (others => '0');
		P_HR_NS210 <= (others => '0');
		P_HR_NS211 <= (others => '0');
		P_HR_NS212 <= (others => '0');
		P_HR_NS213 <= (others => '0');
		P_HR_NS214 <= (others => '0');
		P_HR_NS215 <= (others => '0');
		P_HR_NS216 <= (others => '0');
		P_HR_NS217 <= (others => '0');
		P_HR_NS218 <= (others => '0');
		P_HR_NS219 <= (others => '0');
		P_HR_NS220 <= (others => '0');
		P_HR_NS221 <= (others => '0');
		P_HR_NS222 <= (others => '0');
		P_HR_NS223 <= (others => '0');
		P_HR_NS224 <= (others => '0');
		P_HR_NS225 <= (others => '0');
		P_HR_NS226 <= (others => '0');
		P_HR_NS227 <= (others => '0');
		P_HR_NS228 <= (others => '0');
		P_HR_NS229 <= (others => '0');
		P_HR_NS230 <= (others => '0');
		P_HR_NS231 <= (others => '0');
		P_HR_NS232 <= (others => '0');
		P_HR_NS233 <= (others => '0');
		P_HR_NS234 <= (others => '0');
		P_HR_NS235 <= (others => '0');
		P_HR_NS236 <= (others => '0');
		P_HR_NS237 <= (others => '0');
		P_HR_NS238 <= (others => '0');
		P_HR_NS239 <= (others => '0');
		P_HR_NS240 <= (others => '0');
		P_HR_NS241 <= (others => '0');
		P_HR_NS242 <= (others => '0');
		P_HR_NS243 <= (others => '0');
		P_HR_NS244 <= (others => '0');
		P_HR_NS245 <= (others => '0');
		P_HR_NS246 <= (others => '0');
		P_HR_NS247 <= (others => '0');
		P_HR_NS248 <= (others => '0');
		P_HR_NS249 <= (others => '0');
		P_HR_NS250 <= (others => '0');
		P_HR_NS251 <= (others => '0');
		P_HR_NS252 <= (others => '0');
		P_HR_NS253 <= (others => '0');
		P_HR_NS254 <= (others => '0');
		P_HR_NS255 <= (others => '0');
		P_HR_NS256 <= (others => '0');
		P_HR_NS257 <= (others => '0');
		P_HR_NS258 <= (others => '0');
		P_HR_NS259 <= (others => '0');
		P_HR_NS260 <= (others => '0');
		P_HR_NS261 <= (others => '0');
		P_HR_NS262 <= (others => '0');
		P_HR_NS263 <= (others => '0');
		P_HR_NS264 <= (others => '0');
		P_HR_NS265 <= (others => '0');
		P_HR_NS266 <= (others => '0');
		P_HR_NS267 <= (others => '0');
		P_HR_NS268 <= (others => '0');
		P_HR_NS269 <= (others => '0');
		P_HR_NS270 <= (others => '0');
		P_HR_NS271 <= (others => '0');
		P_HR_NS272 <= (others => '0');
		P_HR_NS273 <= (others => '0');
		P_HR_NS274 <= (others => '0');
		P_HR_NS275 <= (others => '0');
		P_HR_NS276 <= (others => '0');
		P_HR_NS277 <= (others => '0');
		P_HR_NS278 <= (others => '0');
		P_HR_NS279 <= (others => '0');
		P_HR_NS280 <= (others => '0');
		P_HR_NS281 <= (others => '0');
		P_HR_NS282 <= (others => '0');
		P_HR_NS283 <= (others => '0');
		P_HR_NS284 <= (others => '0');
		P_HR_NS285 <= (others => '0');
		P_HR_NS286 <= (others => '0');
		P_HR_NS287 <= (others => '0');
		P_HR_NS288 <= (others => '0');
		P_HR_NS289 <= (others => '0');
		P_HR_NS290 <= (others => '0');
		P_HR_NS291 <= (others => '0');
		P_HR_NS292 <= (others => '0');
		P_HR_NS293 <= (others => '0');
		P_HR_NS294 <= (others => '0');
		P_HR_NS295 <= (others => '0');
		P_HR_NS296 <= (others => '0');
		P_HR_NS297 <= (others => '0');
		P_HR_NS298 <= (others => '0');
		P_HR_NS299 <= (others => '0');
		P_HR_NS300 <= (others => '0');
		P_HR_NS301 <= (others => '0');
		P_HR_NS302 <= (others => '0');
		P_HR_NS303 <= (others => '0');
		P_HR_NS304 <= (others => '0');
		P_HR_NS305 <= (others => '0');
		P_HR_NS306 <= (others => '0');
		P_HR_NS307 <= (others => '0');
		P_HR_NS308 <= (others => '0');
		P_HR_NS309 <= (others => '0');
		P_HR_NS310 <= (others => '0');
		P_HR_NS311 <= (others => '0');
		P_HR_NS312 <= (others => '0');
		P_HR_NS313 <= (others => '0');
		P_HR_NS314 <= (others => '0');
		P_HR_NS315 <= (others => '0');
		P_HR_NS316 <= (others => '0');
		P_HR_NS317 <= (others => '0');
		P_HR_NS318 <= (others => '0');
		P_HR_NS319 <= (others => '0');
		P_HR_NS320 <= (others => '0');
		P_HR_NS321 <= (others => '0');
		P_HR_NS322 <= (others => '0');
		P_HR_NS323 <= (others => '0');
		P_HR_NS324 <= (others => '0');
		P_HR_NS325 <= (others => '0');
		P_HR_NS326 <= (others => '0');
		P_HR_NS327 <= (others => '0');
		P_HR_NS328 <= (others => '0');
		P_HR_NS329 <= (others => '0');
		P_HR_NS330 <= (others => '0');
		P_HR_NS331 <= (others => '0');
		P_HR_NS332 <= (others => '0');
		P_HR_NS333 <= (others => '0');
		P_HR_NS334 <= (others => '0');
		P_HR_NS335 <= (others => '0');
		P_HR_NS336 <= (others => '0');
		P_HR_NS337 <= (others => '0');
		P_HR_NS338 <= (others => '0');
		P_HR_NS339 <= (others => '0');
		P_HR_NS340 <= (others => '0');
		P_HR_NS341 <= (others => '0');
		P_HR_NS342 <= (others => '0');
		P_HR_NS343 <= (others => '0');
		P_HR_NS344 <= (others => '0');
		P_HR_NS345 <= (others => '0');
		P_HR_NS346 <= (others => '0');
		P_HR_NS347 <= (others => '0');
		P_HR_NS348 <= (others => '0');
		P_HR_NS349 <= (others => '0');
		P_HR_NS350 <= (others => '0');
		P_HR_NS351 <= (others => '0');
		P_HR_NS352 <= (others => '0');
		P_HR_NS353 <= (others => '0');
		P_HR_NS354 <= (others => '0');
		P_HR_NS355 <= (others => '0');
		P_HR_NS356 <= (others => '0');
		P_HR_NS357 <= (others => '0');
		P_HR_NS358 <= (others => '0');
		P_HR_NS359 <= (others => '0');
		P_HR_NS360 <= (others => '0');
		P_HR_NS361 <= (others => '0');
		P_HR_NS362 <= (others => '0');
		P_HR_NS363 <= (others => '0');
		P_HR_NS364 <= (others => '0');
		P_HR_NS365 <= (others => '0');
		P_HR_NS366 <= (others => '0');
		P_HR_NS367 <= (others => '0');
		P_HR_NS368 <= (others => '0');
		P_HR_NS369 <= (others => '0');
		P_HR_NS370 <= (others => '0');
		P_HR_NS371 <= (others => '0');
		P_HR_NS372 <= (others => '0');
		P_HR_NS373 <= (others => '0');
		P_HR_NS374 <= (others => '0');
		P_HR_NS375 <= (others => '0');
		P_HR_NS376 <= (others => '0');
		P_HR_NS377 <= (others => '0');
		P_HR_NS378 <= (others => '0');
		P_HR_NS379 <= (others => '0');
		P_HR_NS380 <= (others => '0');
		P_HR_NS381 <= (others => '0');
		P_HR_NS382 <= (others => '0');
		P_HR_NS383 <= (others => '0');
		P_HR_NS384 <= (others => '0');
		P_HR_NS385 <= (others => '0');
		P_HR_NS386 <= (others => '0');
		P_HR_NS387 <= (others => '0');
		P_HR_NS388 <= (others => '0');
		P_HR_NS389 <= (others => '0');
		P_HR_NS390 <= (others => '0');
		P_HR_NS391 <= (others => '0');
		P_HR_NS392 <= (others => '0');
		P_HR_NS393 <= (others => '0');
		P_HR_NS394 <= (others => '0');
		P_HR_NS395 <= (others => '0');
		P_HR_NS396 <= (others => '0');
		P_HR_NS397 <= (others => '0');
		P_HR_NS398 <= (others => '0');
		P_HR_NS399 <= (others => '0');
		P_HR_NS400 <= (others => '0');
		P_HR_NS401 <= (others => '0');
		P_HR_NS402 <= (others => '0');
		P_HR_NS403 <= (others => '0');
		P_HR_NS404 <= (others => '0');
		P_HR_NS405 <= (others => '0');
		P_HR_NS406 <= (others => '0');
		P_HR_NS407 <= (others => '0');
		P_HR_NS408 <= (others => '0');
		P_HR_NS409 <= (others => '0');
		P_HR_NS410 <= (others => '0');
		P_HR_NS411 <= (others => '0');
		P_HR_NS412 <= (others => '0');
		P_HR_NS413 <= (others => '0');
		P_HR_NS414 <= (others => '0');
		P_HR_NS415 <= (others => '0');
		P_HR_NS416 <= (others => '0');
		P_HR_NS417 <= (others => '0');
		P_HR_NS418 <= (others => '0');
		P_HR_NS419 <= (others => '0');
		P_HR_NS420 <= (others => '0');
		P_HR_NS421 <= (others => '0');
		P_HR_NS422 <= (others => '0');
		P_HR_NS423 <= (others => '0');
		P_HR_NS424 <= (others => '0');
		P_HR_NS425 <= (others => '0');
		P_HR_NS426 <= (others => '0');
		P_HR_NS427 <= (others => '0');
		P_HR_NS428 <= (others => '0');
		P_HR_NS429 <= (others => '0');
		P_HR_NS430 <= (others => '0');
		P_HR_NS431 <= (others => '0');
		P_HR_NS432 <= (others => '0');
		P_HR_NS433 <= (others => '0');
		P_HR_NS434 <= (others => '0');
		P_HR_NS435 <= (others => '0');
		P_HR_NS436 <= (others => '0');
		P_HR_NS437 <= (others => '0');
		P_HR_NS438 <= (others => '0');
		P_HR_NS439 <= (others => '0');
		P_HR_NS440 <= (others => '0');
		P_HR_NS441 <= (others => '0');
		P_HR_NS442 <= (others => '0');
		P_HR_NS443 <= (others => '0');
		P_HR_NS444 <= (others => '0');
		P_HR_NS445 <= (others => '0');
		P_HR_NS446 <= (others => '0');
		P_HR_NS447 <= (others => '0');
		P_HR_NS448 <= (others => '0');
		P_HR_NS449 <= (others => '0');
		P_HR_NS450 <= (others => '0');
		P_HR_NS451 <= (others => '0');
		P_HR_NS452 <= (others => '0');
		P_HR_NS453 <= (others => '0');
		P_HR_NS454 <= (others => '0');
		P_HR_NS455 <= (others => '0');
		P_HR_NS456 <= (others => '0');
		P_HR_NS457 <= (others => '0');
		P_HR_NS458 <= (others => '0');	
			
		P_EDA_NS1 <= (others => '0');
		P_EDA_NS2 <= (others => '0');
		P_EDA_NS3 <= (others => '0');
		P_EDA_NS4 <= (others => '0');
		P_EDA_NS5 <= (others => '0');
		P_EDA_NS6 <= (others => '0');
		P_EDA_NS7 <= (others => '0');
		P_EDA_NS8 <= (others => '0');
		P_EDA_NS9 <= (others => '0');
		P_EDA_NS10 <= (others => '0');
		P_EDA_NS11 <= (others => '0');
		P_EDA_NS12 <= (others => '0');
		P_EDA_NS13 <= (others => '0');
		P_EDA_NS14 <= (others => '0');
		P_EDA_NS15 <= (others => '0');
		P_EDA_NS16 <= (others => '0');
		P_EDA_NS17 <= (others => '0');
		P_EDA_NS18 <= (others => '0');
		P_EDA_NS19 <= (others => '0');
		P_EDA_NS20 <= (others => '0');
		P_EDA_NS21 <= (others => '0');
		P_EDA_NS22 <= (others => '0');
		P_EDA_NS23 <= (others => '0');
		P_EDA_NS24 <= (others => '0');
		P_EDA_NS25 <= (others => '0');
		P_EDA_NS26 <= (others => '0');
		P_EDA_NS27 <= (others => '0');
		P_EDA_NS28 <= (others => '0');
		P_EDA_NS29 <= (others => '0');
		P_EDA_NS30 <= (others => '0');
		P_EDA_NS31 <= (others => '0');
		P_EDA_NS32 <= (others => '0');
		P_EDA_NS33 <= (others => '0');
		P_EDA_NS34 <= (others => '0');
		P_EDA_NS35 <= (others => '0');
		P_EDA_NS36 <= (others => '0');
		P_EDA_NS37 <= (others => '0');
		P_EDA_NS38 <= (others => '0');
		P_EDA_NS39 <= (others => '0');
		P_EDA_NS40 <= (others => '0');
		P_EDA_NS41 <= (others => '0');
		P_EDA_NS42 <= (others => '0');
		P_EDA_NS43 <= (others => '0');
		P_EDA_NS44 <= (others => '0');
		P_EDA_NS45 <= (others => '0');
		P_EDA_NS46 <= (others => '0');
		P_EDA_NS47 <= (others => '0');
		P_EDA_NS48 <= (others => '0');
		P_EDA_NS49 <= (others => '0');
		P_EDA_NS50 <= (others => '0');
		P_EDA_NS51 <= (others => '0');
		P_EDA_NS52 <= (others => '0');
		P_EDA_NS53 <= (others => '0');
		P_EDA_NS54 <= (others => '0');
		P_EDA_NS55 <= (others => '0');
		P_EDA_NS56 <= (others => '0');
		P_EDA_NS57 <= (others => '0');
		P_EDA_NS58 <= (others => '0');
		P_EDA_NS59 <= (others => '0');
		P_EDA_NS60 <= (others => '0');
		P_EDA_NS61 <= (others => '0');
		P_EDA_NS62 <= (others => '0');
		P_EDA_NS63 <= (others => '0');
		P_EDA_NS64 <= (others => '0');
		P_EDA_NS65 <= (others => '0');
		P_EDA_NS66 <= (others => '0');
		P_EDA_NS67 <= (others => '0');	

		P_TEMP_NS <= (others => '0');	
		P_EDA_NS <= (others => '0');	
		P_HR_NS <= (others => '0');		
		
		not_stress_score <= (others => '0');		
			
		elsif (rising_edge(clk)) then
		if state = NORMAL then
			case temp is
				when "011100000" => P_TEMP_NS <= "000000000001" + P_TEMP_NS1;
				when "011100001" => P_TEMP_NS <= "000000110101" + P_TEMP_NS2;
				when "011100010" => P_TEMP_NS <= "000011110110" + P_TEMP_NS3;
				when "011100011" => P_TEMP_NS <= "001001111011" + P_TEMP_NS4;
				when "011100100" => P_TEMP_NS <= "001000010000" + P_TEMP_NS5;
				when "011100101" => P_TEMP_NS <= "000010010100" + P_TEMP_NS6;
				when "011100110" => P_TEMP_NS <= "000011000001" + P_TEMP_NS7;
				when "011100111" => P_TEMP_NS <= "000010000001" + P_TEMP_NS8;
				when "011101000" => P_TEMP_NS <= "000000101000" + P_TEMP_NS9;
				when "011101001" => P_TEMP_NS <= "000001000010" + P_TEMP_NS10;
				when "011101010" => P_TEMP_NS <= "000000101010" + P_TEMP_NS11;
				when "011101011" => P_TEMP_NS <= "000000000100" + P_TEMP_NS12;
				when "011101100" => P_TEMP_NS <= "000000000011" + P_TEMP_NS13;
				when "011101101" => P_TEMP_NS <= "000000000011" + P_TEMP_NS14;
				when "011101110" => P_TEMP_NS <= "000000001001" + P_TEMP_NS15;
				when "011101111" => P_TEMP_NS <= "000000001000" + P_TEMP_NS16;
				when "011110000" => P_TEMP_NS <= "000000001000" + P_TEMP_NS17;
				when "011110001" => P_TEMP_NS <= "000000001000" + P_TEMP_NS18;
				when "011110010" => P_TEMP_NS <= "000000001000" + P_TEMP_NS19;
				when "011110011" => P_TEMP_NS <= "000000000111" + P_TEMP_NS20;
				when "011110100" => P_TEMP_NS <= "000000000111" + P_TEMP_NS21;
				when "011110101" => P_TEMP_NS <= "000000000111" + P_TEMP_NS22;
				when "011110110" => P_TEMP_NS <= "000001100000" + P_TEMP_NS23;
				when "011110111" => P_TEMP_NS <= "000110100010" + P_TEMP_NS24;
				when "011111000" => P_TEMP_NS <= "000101001111" + P_TEMP_NS25;
				when "011111001" => P_TEMP_NS <= "000010001010" + P_TEMP_NS26;
				when "011111010" => P_TEMP_NS <= "000100101011" + P_TEMP_NS27;
				when "011111011" => P_TEMP_NS <= "001110100000" + P_TEMP_NS28;
				when "011111100" => P_TEMP_NS <= "000100101110" + P_TEMP_NS29;
				when "011111101" => P_TEMP_NS <= "000110111000" + P_TEMP_NS30;
				when "011111110" => P_TEMP_NS <= "000011101101" + P_TEMP_NS31;
				when "011111111" => P_TEMP_NS <= "000100011000" + P_TEMP_NS32;
				when "100000000" => P_TEMP_NS <= "001001010110" + P_TEMP_NS33;
				when "100000001" => P_TEMP_NS <= "001000010000" + P_TEMP_NS34;
				when "100000010" => P_TEMP_NS <= "000010010111" + P_TEMP_NS35;
				when "100000011" => P_TEMP_NS <= "000001101011" + P_TEMP_NS36;
				when "100000100" => P_TEMP_NS <= "000010001010" + P_TEMP_NS37;
				when "100000101" => P_TEMP_NS <= "000001111001" + P_TEMP_NS38;
				when "100000110" => P_TEMP_NS <= "000001101010" + P_TEMP_NS39;
				when "100000111" => P_TEMP_NS <= "000100110011" + P_TEMP_NS40;
				when "100001000" => P_TEMP_NS <= "001000100001" + P_TEMP_NS41;
				when "100001001" => P_TEMP_NS <= "001011000100" + P_TEMP_NS42;
				when "100001010" => P_TEMP_NS <= "000111000000" + P_TEMP_NS43;
				when "100001011" => P_TEMP_NS <= "001000001101" + P_TEMP_NS44;
				when "100001100" => P_TEMP_NS <= "000000001100" + P_TEMP_NS45;
				when "100001101" => P_TEMP_NS <= "000000001001" + P_TEMP_NS46;
				when "100001110" => P_TEMP_NS <= "000000001010" + P_TEMP_NS47;
				when "100001111" => P_TEMP_NS <= "000000001100" + P_TEMP_NS48;
				when "100010000" => P_TEMP_NS <= "000000001111" + P_TEMP_NS49;
				when "100010001" => P_TEMP_NS <= "000000010011" + P_TEMP_NS50;
				when "100010010" => P_TEMP_NS <= "000000001100" + P_TEMP_NS51;
				when "100010011" => P_TEMP_NS <= "000000000010" + P_TEMP_NS52;
				when  others     => P_TEMP_NS <= "000000000001";
			end case;	
		
        case hr is
				when "00000000001" => P_HR_NS <= "000000000100" + P_HR_NS1;
				when "00000000011" => P_HR_NS <= "000000000100" + P_HR_NS2;
				when "00000000100" => P_HR_NS <= "000000000100" + P_HR_NS3;
				when "00000000111" => P_HR_NS <= "000000000100" + P_HR_NS4;
				when "00000001000" => P_HR_NS <= "000000000100" + P_HR_NS5;
				when "00000001001" => P_HR_NS <= "000000001011" + P_HR_NS6;
				when "00000001010" => P_HR_NS <= "000000000100" + P_HR_NS7;
				when "00000001101" => P_HR_NS <= "000000000111" + P_HR_NS8;
				when "00000001110" => P_HR_NS <= "000000000100" + P_HR_NS9;
				when "00000010000" => P_HR_NS <= "000000000100" + P_HR_NS10;
				when "00000010001" => P_HR_NS <= "000000001011" + P_HR_NS11;
				when "00000010011" => P_HR_NS <= "000000000100" + P_HR_NS12;
				when "00000010101" => P_HR_NS <= "000000000100" + P_HR_NS13;
				when "00000011100" => P_HR_NS <= "000000001011" + P_HR_NS14;
				when "00000011101" => P_HR_NS <= "000000000100" + P_HR_NS15;
				when "00000101001" => P_HR_NS <= "000000000100" + P_HR_NS16;
				when "00000110101" => P_HR_NS <= "000000000100" + P_HR_NS17;
				when "00000111000" => P_HR_NS <= "000000000100" + P_HR_NS18;
				when "00001000001" => P_HR_NS <= "000000000100" + P_HR_NS19;
				when "00001001100" => P_HR_NS <= "000000000100" + P_HR_NS20;
				when "00001010011" => P_HR_NS <= "000000000111" + P_HR_NS21;
				when "00001011100" => P_HR_NS <= "000000000100" + P_HR_NS22;
				when "00001101001" => P_HR_NS <= "000000000100" + P_HR_NS23;
				when "00001101100" => P_HR_NS <= "000000000100" + P_HR_NS24;
				when "00001101111" => P_HR_NS <= "000000000100" + P_HR_NS25;
				when "00001110000" => P_HR_NS <= "000000000100" + P_HR_NS26;
				when "00001110101" => P_HR_NS <= "000000000100" + P_HR_NS27;
				when "00001110110" => P_HR_NS <= "000000000100" + P_HR_NS28;
				when "00001111000" => P_HR_NS <= "000000000100" + P_HR_NS29;
				when "00001111110" => P_HR_NS <= "000000000100" + P_HR_NS30;
				when "00001111111" => P_HR_NS <= "000000000100" + P_HR_NS31;
				when "00010000000" => P_HR_NS <= "000000000100" + P_HR_NS32;
				when "00010000010" => P_HR_NS <= "000000000100" + P_HR_NS33;
				when "00010000100" => P_HR_NS <= "000000000100" + P_HR_NS34;
				when "00010000101" => P_HR_NS <= "000000000100" + P_HR_NS35;
				when "00010000110" => P_HR_NS <= "000000000100" + P_HR_NS36;
				when "00010001010" => P_HR_NS <= "000000000111" + P_HR_NS37;
				when "00010001011" => P_HR_NS <= "000000000111" + P_HR_NS38;
				when "00010001100" => P_HR_NS <= "000000000100" + P_HR_NS39;
				when "00010010010" => P_HR_NS <= "000000000100" + P_HR_NS40;
				when "00010010100" => P_HR_NS <= "000000000100" + P_HR_NS41;
				when "00010011100" => P_HR_NS <= "000000000100" + P_HR_NS42;
				when "00010100001" => P_HR_NS <= "000000000100" + P_HR_NS43;
				when "00010100101" => P_HR_NS <= "000000001011" + P_HR_NS44;
				when "00010100110" => P_HR_NS <= "000000000100" + P_HR_NS45;
				when "00010100111" => P_HR_NS <= "000000000111" + P_HR_NS46;
				when "00010101001" => P_HR_NS <= "000000001011" + P_HR_NS47;
				when "00010101010" => P_HR_NS <= "000000000100" + P_HR_NS48;
				when "00010101011" => P_HR_NS <= "000000001011" + P_HR_NS49;
				when "00010101101" => P_HR_NS <= "000000001011" + P_HR_NS50;
				when "00010101110" => P_HR_NS <= "000000001011" + P_HR_NS51;
				when "00010101111" => P_HR_NS <= "000000010101" + P_HR_NS52;
				when "00010110000" => P_HR_NS <= "000000010101" + P_HR_NS53;
				when "00010110001" => P_HR_NS <= "000000010010" + P_HR_NS54;
				when "00010110010" => P_HR_NS <= "000000000111" + P_HR_NS55;
				when "00010110011" => P_HR_NS <= "000000100111" + P_HR_NS56;
				when "00010110100" => P_HR_NS <= "000000001110" + P_HR_NS57;
				when "00010110101" => P_HR_NS <= "000000000111" + P_HR_NS58;
				when "00010110110" => P_HR_NS <= "000000000111" + P_HR_NS59;
				when "00010110111" => P_HR_NS <= "000000001011" + P_HR_NS60;
				when "00010111000" => P_HR_NS <= "000000001011" + P_HR_NS61;
				when "00010111001" => P_HR_NS <= "000000010010" + P_HR_NS62;
				when "00010111010" => P_HR_NS <= "000000001110" + P_HR_NS63;
				when "00010111011" => P_HR_NS <= "000000001011" + P_HR_NS64;
				when "00010111100" => P_HR_NS <= "000000000111" + P_HR_NS65;
				when "00010111101" => P_HR_NS <= "000000000100" + P_HR_NS66;
				when "00010111110" => P_HR_NS <= "000000001011" + P_HR_NS67;
				when "00010111111" => P_HR_NS <= "000000001011" + P_HR_NS68;
				when "00011000000" => P_HR_NS <= "000000000100" + P_HR_NS69;
				when "00011000010" => P_HR_NS <= "000000000100" + P_HR_NS70;
				when "00011000011" => P_HR_NS <= "000000000100" + P_HR_NS71;
				when "00011000100" => P_HR_NS <= "000000001011" + P_HR_NS72;
				when "00011000101" => P_HR_NS <= "000000000111" + P_HR_NS73;
				when "00011100010" => P_HR_NS <= "000000000100" + P_HR_NS74;
				when "00011100011" => P_HR_NS <= "000000000100" + P_HR_NS75;
				when "00011100101" => P_HR_NS <= "000000000100" + P_HR_NS76;
				when "00011100110" => P_HR_NS <= "000000000100" + P_HR_NS77;
				when "00011101001" => P_HR_NS <= "000000000100" + P_HR_NS78;
				when "00011101010" => P_HR_NS <= "000000000100" + P_HR_NS79;
				when "00011101011" => P_HR_NS <= "000000000111" + P_HR_NS80;
				when "00011101101" => P_HR_NS <= "000000000100" + P_HR_NS81;
				when "00011101111" => P_HR_NS <= "000000000100" + P_HR_NS82;
				when "00011110000" => P_HR_NS <= "000000001011" + P_HR_NS83;
				when "00011110011" => P_HR_NS <= "000000000100" + P_HR_NS84;
				when "00011110101" => P_HR_NS <= "000000000111" + P_HR_NS85;
				when "00011110110" => P_HR_NS <= "000000000100" + P_HR_NS86;
				when "00011111000" => P_HR_NS <= "000000000111" + P_HR_NS87;
				when "00011111001" => P_HR_NS <= "000000001011" + P_HR_NS88;
				when "00011111010" => P_HR_NS <= "000000000100" + P_HR_NS89;
				when "00011111011" => P_HR_NS <= "000000000100" + P_HR_NS90;
				when "00011111100" => P_HR_NS <= "000000000100" + P_HR_NS91;
				when "00011111101" => P_HR_NS <= "000000000100" + P_HR_NS92;
				when "00011111110" => P_HR_NS <= "000000000111" + P_HR_NS93;
				when "00011111111" => P_HR_NS <= "000000000100" + P_HR_NS94;
				when "00100000000" => P_HR_NS <= "000000001110" + P_HR_NS95;
				when "00100000001" => P_HR_NS <= "000000001110" + P_HR_NS96;
				when "00100000010" => P_HR_NS <= "000000000111" + P_HR_NS97;
				when "00100000011" => P_HR_NS <= "000000001011" + P_HR_NS98;
				when "00100000100" => P_HR_NS <= "000000001011" + P_HR_NS99;
				when "00100000101" => P_HR_NS <= "000000000100" + P_HR_NS100;
				when "00100000110" => P_HR_NS <= "000000001011" + P_HR_NS101;
				when "00100000111" => P_HR_NS <= "000000000111" + P_HR_NS102;
				when "00100001000" => P_HR_NS <= "000000000100" + P_HR_NS103;
				when "00100001001" => P_HR_NS <= "000000000111" + P_HR_NS104;
				when "00100001010" => P_HR_NS <= "000000001011" + P_HR_NS105;
				when "00100001011" => P_HR_NS <= "000000001011" + P_HR_NS106;
				when "00100001100" => P_HR_NS <= "000000001110" + P_HR_NS107;
				when "00100001101" => P_HR_NS <= "000000001110" + P_HR_NS108;
				when "00100001110" => P_HR_NS <= "000000000111" + P_HR_NS109;
				when "00100001111" => P_HR_NS <= "000000010101" + P_HR_NS110;
				when "00100010000" => P_HR_NS <= "000000001110" + P_HR_NS111;
				when "00100010011" => P_HR_NS <= "000000000111" + P_HR_NS112;
				when "00100010100" => P_HR_NS <= "000000000100" + P_HR_NS113;
				when "00100010110" => P_HR_NS <= "000000000100" + P_HR_NS114;
				when "00100010111" => P_HR_NS <= "000000000100" + P_HR_NS115;
				when "00100011000" => P_HR_NS <= "000000001011" + P_HR_NS116;
				when "00100011001" => P_HR_NS <= "000000000111" + P_HR_NS117;
				when "00100011010" => P_HR_NS <= "000000000100" + P_HR_NS118;
				when "00100011011" => P_HR_NS <= "000000000100" + P_HR_NS119;
				when "00100011100" => P_HR_NS <= "000000000111" + P_HR_NS120;
				when "00100011110" => P_HR_NS <= "000000000111" + P_HR_NS121;
				when "00100011111" => P_HR_NS <= "000000000100" + P_HR_NS122;
				when "00100100000" => P_HR_NS <= "000000000111" + P_HR_NS123;
				when "00100100001" => P_HR_NS <= "000000001011" + P_HR_NS124;
				when "00100100010" => P_HR_NS <= "000000000100" + P_HR_NS125;
				when "00100100011" => P_HR_NS <= "000000000100" + P_HR_NS126;
				when "00100100100" => P_HR_NS <= "000000000100" + P_HR_NS127;
				when "00100100110" => P_HR_NS <= "000000000100" + P_HR_NS128;
				when "00100101001" => P_HR_NS <= "000000001011" + P_HR_NS129;
				when "00100101010" => P_HR_NS <= "000000000111" + P_HR_NS130;
				when "00100101011" => P_HR_NS <= "000000001011" + P_HR_NS131;
				when "00100101100" => P_HR_NS <= "000000000100" + P_HR_NS132;
				when "00100101101" => P_HR_NS <= "000000000111" + P_HR_NS133;
				when "00100101110" => P_HR_NS <= "000000000100" + P_HR_NS134;
				when "00100110000" => P_HR_NS <= "000000000100" + P_HR_NS135;
				when "00100110010" => P_HR_NS <= "000000000111" + P_HR_NS136;
				when "00100110011" => P_HR_NS <= "000000000111" + P_HR_NS137;
				when "00100110100" => P_HR_NS <= "000000000100" + P_HR_NS138;
				when "00100110110" => P_HR_NS <= "000000000111" + P_HR_NS139;
				when "00100111000" => P_HR_NS <= "000000000100" + P_HR_NS140;
				when "00100111010" => P_HR_NS <= "000000000100" + P_HR_NS141;
				when "00100111011" => P_HR_NS <= "000000001011" + P_HR_NS142;
				when "00100111100" => P_HR_NS <= "000000000100" + P_HR_NS143;
				when "00100111110" => P_HR_NS <= "000000000111" + P_HR_NS144;
				when "00100111111" => P_HR_NS <= "000000000100" + P_HR_NS145;
				when "00101000000" => P_HR_NS <= "000000001011" + P_HR_NS146;
				when "00101000010" => P_HR_NS <= "000000000111" + P_HR_NS147;
				when "00101000011" => P_HR_NS <= "000000000111" + P_HR_NS148;
				when "00101000100" => P_HR_NS <= "000000000100" + P_HR_NS149;
				when "00101000101" => P_HR_NS <= "000000000100" + P_HR_NS150;
				when "00101000110" => P_HR_NS <= "000000000111" + P_HR_NS151;
				when "00101000111" => P_HR_NS <= "000000000111" + P_HR_NS152;
				when "00101001000" => P_HR_NS <= "000000000111" + P_HR_NS153;
				when "00101001011" => P_HR_NS <= "000000001011" + P_HR_NS154;
				when "00101001110" => P_HR_NS <= "000000000100" + P_HR_NS155;
				when "00101001111" => P_HR_NS <= "000000000111" + P_HR_NS156;
				when "00101010000" => P_HR_NS <= "000000000100" + P_HR_NS157;
				when "00101010001" => P_HR_NS <= "000000001110" + P_HR_NS158;
				when "00101010010" => P_HR_NS <= "000000001110" + P_HR_NS159;
				when "00101010100" => P_HR_NS <= "000000010101" + P_HR_NS160;
				when "00101010101" => P_HR_NS <= "000000000111" + P_HR_NS161;
				when "00101010110" => P_HR_NS <= "000000000111" + P_HR_NS162;
				when "00101010111" => P_HR_NS <= "000000001110" + P_HR_NS163;
				when "00101011000" => P_HR_NS <= "000000010010" + P_HR_NS164;
				when "00101011001" => P_HR_NS <= "000000000111" + P_HR_NS165;
				when "00101011010" => P_HR_NS <= "000000010010" + P_HR_NS166;
				when "00101011011" => P_HR_NS <= "000000001110" + P_HR_NS167;
				when "00101011100" => P_HR_NS <= "000000000111" + P_HR_NS168;
				when "00101011101" => P_HR_NS <= "000000010101" + P_HR_NS169;
				when "00101011110" => P_HR_NS <= "000000001011" + P_HR_NS170;
				when "00101011111" => P_HR_NS <= "000000000100" + P_HR_NS171;
				when "00101100000" => P_HR_NS <= "000000000111" + P_HR_NS172;
				when "00101100001" => P_HR_NS <= "000000001110" + P_HR_NS173;
				when "00101100010" => P_HR_NS <= "000000010010" + P_HR_NS174;
				when "00101100011" => P_HR_NS <= "000000001110" + P_HR_NS175;
				when "00101100100" => P_HR_NS <= "000000010010" + P_HR_NS176;
				when "00101100101" => P_HR_NS <= "000000011001" + P_HR_NS177;
				when "00101100110" => P_HR_NS <= "000000000100" + P_HR_NS178;
				when "00101100111" => P_HR_NS <= "000000100011" + P_HR_NS179;
				when "00101101000" => P_HR_NS <= "000000010101" + P_HR_NS180;
				when "00101101001" => P_HR_NS <= "000000100011" + P_HR_NS181;
				when "00101101010" => P_HR_NS <= "000000100111" + P_HR_NS182;
				when "00101101011" => P_HR_NS <= "000000011001" + P_HR_NS183;
				when "00101101100" => P_HR_NS <= "000000011001" + P_HR_NS184;
				when "00101101101" => P_HR_NS <= "000000011100" + P_HR_NS185;
				when "00101101110" => P_HR_NS <= "000000111100" + P_HR_NS186;
				when "00101101111" => P_HR_NS <= "000000100011" + P_HR_NS187;
				when "00101110000" => P_HR_NS <= "000000110001" + P_HR_NS188;
				when "00101110001" => P_HR_NS <= "000000011001" + P_HR_NS189;
				when "00101110010" => P_HR_NS <= "000000111100" + P_HR_NS190;
				when "00101110011" => P_HR_NS <= "000000100000" + P_HR_NS191;
				when "00101110100" => P_HR_NS <= "000000010101" + P_HR_NS192;
				when "00101110101" => P_HR_NS <= "000000011100" + P_HR_NS193;
				when "00101110110" => P_HR_NS <= "000000011100" + P_HR_NS194;
				when "00101110111" => P_HR_NS <= "000000111100" + P_HR_NS195;
				when "00101111000" => P_HR_NS <= "000000111000" + P_HR_NS196;
				when "00101111001" => P_HR_NS <= "000000100011" + P_HR_NS197;
				when "00101111010" => P_HR_NS <= "000000100111" + P_HR_NS198;
				when "00101111011" => P_HR_NS <= "000000100000" + P_HR_NS199;
				when "00101111100" => P_HR_NS <= "000000010101" + P_HR_NS200;
				when "00101111101" => P_HR_NS <= "000001000110" + P_HR_NS201;
				when "00101111110" => P_HR_NS <= "000000100111" + P_HR_NS202;
				when "00101111111" => P_HR_NS <= "000000010010" + P_HR_NS203;
				when "00110000000" => P_HR_NS <= "000001000011" + P_HR_NS204;
				when "00110000001" => P_HR_NS <= "000000011100" + P_HR_NS205;
				when "00110000010" => P_HR_NS <= "000000010101" + P_HR_NS206;
				when "00110000011" => P_HR_NS <= "000000110101" + P_HR_NS207;
				when "00110000100" => P_HR_NS <= "000001011000" + P_HR_NS208;
				when "00110000101" => P_HR_NS <= "000000100011" + P_HR_NS209;
				when "00110000110" => P_HR_NS <= "000000110101" + P_HR_NS210;
				when "00110000111" => P_HR_NS <= "000000111100" + P_HR_NS211;
				when "00110001000" => P_HR_NS <= "000000100111" + P_HR_NS212;
				when "00110001001" => P_HR_NS <= "000001101101" + P_HR_NS213;
				when "00110001010" => P_HR_NS <= "000000110001" + P_HR_NS214;
				when "00110001011" => P_HR_NS <= "000000110101" + P_HR_NS215;
				when "00110001100" => P_HR_NS <= "000001000110" + P_HR_NS216;
				when "00110001101" => P_HR_NS <= "000000110001" + P_HR_NS217;
				when "00110001110" => P_HR_NS <= "000001001010" + P_HR_NS218;
				when "00110001111" => P_HR_NS <= "000000100011" + P_HR_NS219;
				when "00110010000" => P_HR_NS <= "000001110001" + P_HR_NS220;
				when "00110010001" => P_HR_NS <= "000001000110" + P_HR_NS221;
				when "00110010010" => P_HR_NS <= "000001010001" + P_HR_NS222;
				when "00110010011" => P_HR_NS <= "000001001101" + P_HR_NS223;
				when "00110010100" => P_HR_NS <= "000000111100" + P_HR_NS224;
				when "00110010101" => P_HR_NS <= "000001000011" + P_HR_NS225;
				when "00110010110" => P_HR_NS <= "000001000011" + P_HR_NS226;
				when "00110010111" => P_HR_NS <= "000001100011" + P_HR_NS227;
				when "00110011000" => P_HR_NS <= "000001001101" + P_HR_NS228;
				when "00110011001" => P_HR_NS <= "000001001101" + P_HR_NS229;
				when "00110011010" => P_HR_NS <= "000001011100" + P_HR_NS230;
				when "00110011011" => P_HR_NS <= "000000110001" + P_HR_NS231;
				when "00110011100" => P_HR_NS <= "000000111111" + P_HR_NS232;
				when "00110011101" => P_HR_NS <= "000000110001" + P_HR_NS233;
				when "00110011110" => P_HR_NS <= "000000111111" + P_HR_NS234;
				when "00110011111" => P_HR_NS <= "000000101110" + P_HR_NS235;
				when "00110100000" => P_HR_NS <= "000001000110" + P_HR_NS236;
				when "00110100001" => P_HR_NS <= "000001000011" + P_HR_NS237;
				when "00110100010" => P_HR_NS <= "000000111111" + P_HR_NS238;
				when "00110100011" => P_HR_NS <= "000000101010" + P_HR_NS239;
				when "00110100100" => P_HR_NS <= "000000100011" + P_HR_NS240;
				when "00110100101" => P_HR_NS <= "000000111100" + P_HR_NS241;
				when "00110100110" => P_HR_NS <= "000001000011" + P_HR_NS242;
				when "00110100111" => P_HR_NS <= "000000110101" + P_HR_NS243;
				when "00110101000" => P_HR_NS <= "000000110001" + P_HR_NS244;
				when "00110101001" => P_HR_NS <= "000000110101" + P_HR_NS245;
				when "00110101010" => P_HR_NS <= "000001010001" + P_HR_NS246;
				when "00110101011" => P_HR_NS <= "000000101110" + P_HR_NS247;
				when "00110101100" => P_HR_NS <= "000000101010" + P_HR_NS248;
				when "00110101101" => P_HR_NS <= "000001001010" + P_HR_NS249;
				when "00110101110" => P_HR_NS <= "000000100111" + P_HR_NS250;
				when "00110101111" => P_HR_NS <= "000000100011" + P_HR_NS251;
				when "00110110000" => P_HR_NS <= "000001000110" + P_HR_NS252;
				when "00110110001" => P_HR_NS <= "000000010101" + P_HR_NS253;
				when "00110110010" => P_HR_NS <= "000001000011" + P_HR_NS254;
				when "00110110011" => P_HR_NS <= "000000111000" + P_HR_NS255;
				when "00110110100" => P_HR_NS <= "000001010001" + P_HR_NS256;
				when "00110110101" => P_HR_NS <= "000000101010" + P_HR_NS257;
				when "00110110110" => P_HR_NS <= "000000101110" + P_HR_NS258;
				when "00110110111" => P_HR_NS <= "000000101110" + P_HR_NS259;
				when "00110111000" => P_HR_NS <= "000000111000" + P_HR_NS260;
				when "00110111001" => P_HR_NS <= "000000011001" + P_HR_NS261;
				when "00110111010" => P_HR_NS <= "000000110001" + P_HR_NS262;
				when "00110111011" => P_HR_NS <= "000001000110" + P_HR_NS263;
				when "00110111100" => P_HR_NS <= "000000110001" + P_HR_NS264;
				when "00110111101" => P_HR_NS <= "000000100000" + P_HR_NS265;
				when "00110111110" => P_HR_NS <= "000000101010" + P_HR_NS266;
				when "00110111111" => P_HR_NS <= "000000110101" + P_HR_NS267;
				when "00111000000" => P_HR_NS <= "000000100111" + P_HR_NS268;
				when "00111000001" => P_HR_NS <= "000000111100" + P_HR_NS269;
				when "00111000010" => P_HR_NS <= "000001000110" + P_HR_NS270;
				when "00111000011" => P_HR_NS <= "000000010010" + P_HR_NS271;
				when "00111000100" => P_HR_NS <= "000000100011" + P_HR_NS272;
				when "00111000101" => P_HR_NS <= "000000101110" + P_HR_NS273;
				when "00111000110" => P_HR_NS <= "000000011100" + P_HR_NS274;
				when "00111000111" => P_HR_NS <= "000000011001" + P_HR_NS275;
				when "00111001000" => P_HR_NS <= "000000010101" + P_HR_NS276;
				when "00111001001" => P_HR_NS <= "000000111000" + P_HR_NS277;
				when "00111001010" => P_HR_NS <= "000000110001" + P_HR_NS278;
				when "00111001011" => P_HR_NS <= "000000010010" + P_HR_NS279;
				when "00111001100" => P_HR_NS <= "000000100111" + P_HR_NS280;
				when "00111001101" => P_HR_NS <= "000000010101" + P_HR_NS281;
				when "00111001110" => P_HR_NS <= "000000101010" + P_HR_NS282;
				when "00111001111" => P_HR_NS <= "000000110001" + P_HR_NS283;
				when "00111010000" => P_HR_NS <= "000000000111" + P_HR_NS284;
				when "00111010001" => P_HR_NS <= "000000011100" + P_HR_NS285;
				when "00111010010" => P_HR_NS <= "000000011100" + P_HR_NS286;
				when "00111010011" => P_HR_NS <= "000001000011" + P_HR_NS287;
				when "00111010100" => P_HR_NS <= "000000100000" + P_HR_NS288;
				when "00111010101" => P_HR_NS <= "000000110001" + P_HR_NS289;
				when "00111010110" => P_HR_NS <= "000000011100" + P_HR_NS290;
				when "00111010111" => P_HR_NS <= "000000111000" + P_HR_NS291;
				when "00111011000" => P_HR_NS <= "000000100011" + P_HR_NS292;
				when "00111011001" => P_HR_NS <= "000001000110" + P_HR_NS293;
				when "00111011010" => P_HR_NS <= "000000011100" + P_HR_NS294;
				when "00111011011" => P_HR_NS <= "000000100000" + P_HR_NS295;
				when "00111011100" => P_HR_NS <= "000000100111" + P_HR_NS296;
				when "00111011101" => P_HR_NS <= "000000110001" + P_HR_NS297;
				when "00111011110" => P_HR_NS <= "000000011100" + P_HR_NS298;
				when "00111011111" => P_HR_NS <= "000001001101" + P_HR_NS299;
				when "00111100000" => P_HR_NS <= "000000011100" + P_HR_NS300;
				when "00111100001" => P_HR_NS <= "000000101110" + P_HR_NS301;
				when "00111100010" => P_HR_NS <= "000000001011" + P_HR_NS302;
				when "00111100011" => P_HR_NS <= "000000100111" + P_HR_NS303;
				when "00111100100" => P_HR_NS <= "000000001011" + P_HR_NS304;
				when "00111100101" => P_HR_NS <= "000000100111" + P_HR_NS305;
				when "00111100110" => P_HR_NS <= "000001000110" + P_HR_NS306;
				when "00111100111" => P_HR_NS <= "000000010101" + P_HR_NS307;
				when "00111101000" => P_HR_NS <= "000000011100" + P_HR_NS308;
				when "00111101001" => P_HR_NS <= "000000010010" + P_HR_NS309;
				when "00111101010" => P_HR_NS <= "000000010101" + P_HR_NS310;
				when "00111101011" => P_HR_NS <= "000000101110" + P_HR_NS311;
				when "00111101100" => P_HR_NS <= "000000010101" + P_HR_NS312;
				when "00111101101" => P_HR_NS <= "000000100000" + P_HR_NS313;
				when "00111101110" => P_HR_NS <= "000000000111" + P_HR_NS314;
				when "00111101111" => P_HR_NS <= "000000100011" + P_HR_NS315;
				when "00111110000" => P_HR_NS <= "000000110101" + P_HR_NS316;
				when "00111110001" => P_HR_NS <= "000000010010" + P_HR_NS317;
				when "00111110010" => P_HR_NS <= "000000010101" + P_HR_NS318;
				when "00111110011" => P_HR_NS <= "000000111100" + P_HR_NS319;
				when "00111110100" => P_HR_NS <= "000000011001" + P_HR_NS320;
				when "00111110101" => P_HR_NS <= "000000010010" + P_HR_NS321;
				when "00111110110" => P_HR_NS <= "000000001110" + P_HR_NS322;
				when "00111110111" => P_HR_NS <= "000000110001" + P_HR_NS323;
				when "00111111000" => P_HR_NS <= "000000001110" + P_HR_NS324;
				when "00111111001" => P_HR_NS <= "000000101110" + P_HR_NS325;
				when "00111111010" => P_HR_NS <= "000000001011" + P_HR_NS326;
				when "00111111011" => P_HR_NS <= "000000011001" + P_HR_NS327;
				when "00111111100" => P_HR_NS <= "000000100011" + P_HR_NS328;
				when "00111111101" => P_HR_NS <= "000000010010" + P_HR_NS329;
				when "00111111110" => P_HR_NS <= "000000010101" + P_HR_NS330;
				when "00111111111" => P_HR_NS <= "000000100111" + P_HR_NS331;
				when "01000000000" => P_HR_NS <= "000000011001" + P_HR_NS332;
				when "01000000001" => P_HR_NS <= "000000000111" + P_HR_NS333;
				when "01000000010" => P_HR_NS <= "000000011001" + P_HR_NS334;
				when "01000000011" => P_HR_NS <= "000000110001" + P_HR_NS335;
				when "01000000100" => P_HR_NS <= "000000011100" + P_HR_NS336;
				when "01000000101" => P_HR_NS <= "000000001110" + P_HR_NS337;
				when "01000000110" => P_HR_NS <= "000000011001" + P_HR_NS338;
				when "01000000111" => P_HR_NS <= "000000111100" + P_HR_NS339;
				when "01000001000" => P_HR_NS <= "000000011100" + P_HR_NS340;
				when "01000001001" => P_HR_NS <= "000000011100" + P_HR_NS341;
				when "01000001010" => P_HR_NS <= "000000010010" + P_HR_NS342;
				when "01000001011" => P_HR_NS <= "000000110101" + P_HR_NS343;
				when "01000001100" => P_HR_NS <= "000000011001" + P_HR_NS344;
				when "01000001101" => P_HR_NS <= "000000001011" + P_HR_NS345;
				when "01000001110" => P_HR_NS <= "000000010101" + P_HR_NS346;
				when "01000001111" => P_HR_NS <= "000000101110" + P_HR_NS347;
				when "01000010000" => P_HR_NS <= "000000100000" + P_HR_NS348;
				when "01000010001" => P_HR_NS <= "000000010101" + P_HR_NS349;
				when "01000010010" => P_HR_NS <= "000000011001" + P_HR_NS350;
				when "01000010011" => P_HR_NS <= "000000011100" + P_HR_NS351;
				when "01000010100" => P_HR_NS <= "000000111000" + P_HR_NS352;
				when "01000010101" => P_HR_NS <= "000000010010" + P_HR_NS353;
				when "01000010110" => P_HR_NS <= "000000011100" + P_HR_NS354;
				when "01000010111" => P_HR_NS <= "000000010010" + P_HR_NS355;
				when "01000011000" => P_HR_NS <= "000000100000" + P_HR_NS356;
				when "01000011001" => P_HR_NS <= "000000001110" + P_HR_NS357;
				when "01000011010" => P_HR_NS <= "000000101010" + P_HR_NS358;
				when "01000011011" => P_HR_NS <= "000000001110" + P_HR_NS359;
				when "01000011100" => P_HR_NS <= "000000100011" + P_HR_NS360;
				when "01000011101" => P_HR_NS <= "000000010101" + P_HR_NS361;
				when "01000011110" => P_HR_NS <= "000000001110" + P_HR_NS362;
				when "01000011111" => P_HR_NS <= "000000011001" + P_HR_NS363;
				when "01000100000" => P_HR_NS <= "000000100000" + P_HR_NS364;
				when "01000100001" => P_HR_NS <= "000000011001" + P_HR_NS365;
				when "01000100010" => P_HR_NS <= "000000010010" + P_HR_NS366;
				when "01000100011" => P_HR_NS <= "000000001110" + P_HR_NS367;
				when "01000100100" => P_HR_NS <= "000000010101" + P_HR_NS368;
				when "01000100101" => P_HR_NS <= "000000010010" + P_HR_NS369;
				when "01000100110" => P_HR_NS <= "000000011100" + P_HR_NS370;
				when "01000100111" => P_HR_NS <= "000000011001" + P_HR_NS371;
				when "01000101000" => P_HR_NS <= "000000010010" + P_HR_NS372;
				when "01000101001" => P_HR_NS <= "000000000100" + P_HR_NS373;
				when "01000101010" => P_HR_NS <= "000000100111" + P_HR_NS374;
				when "01000101011" => P_HR_NS <= "000000011001" + P_HR_NS375;
				when "01000101100" => P_HR_NS <= "000000001011" + P_HR_NS376;
				when "01000101101" => P_HR_NS <= "000000001011" + P_HR_NS377;
				when "01000101110" => P_HR_NS <= "000000100011" + P_HR_NS378;
				when "01000101111" => P_HR_NS <= "000000001110" + P_HR_NS379;
				when "01000110000" => P_HR_NS <= "000000000111" + P_HR_NS380;
				when "01000110001" => P_HR_NS <= "000000010101" + P_HR_NS381;
				when "01000110010" => P_HR_NS <= "000000001110" + P_HR_NS382;
				when "01000110011" => P_HR_NS <= "000000000100" + P_HR_NS383;
				when "01000110100" => P_HR_NS <= "000000010010" + P_HR_NS384;
				when "01000110110" => P_HR_NS <= "000000001110" + P_HR_NS385;
				when "01000110111" => P_HR_NS <= "000000000111" + P_HR_NS386;
				when "01000111000" => P_HR_NS <= "000000001110" + P_HR_NS387;
				when "01000111001" => P_HR_NS <= "000000100000" + P_HR_NS388;
				when "01000111010" => P_HR_NS <= "000000000100" + P_HR_NS389;
				when "01000111011" => P_HR_NS <= "000000001110" + P_HR_NS390;
				when "01000111100" => P_HR_NS <= "000000010101" + P_HR_NS391;
				when "01000111101" => P_HR_NS <= "000000001011" + P_HR_NS392;
				when "01000111110" => P_HR_NS <= "000000001011" + P_HR_NS393;
				when "01000111111" => P_HR_NS <= "000000001110" + P_HR_NS394;
				when "01001000000" => P_HR_NS <= "000000001011" + P_HR_NS395;
				when "01001000001" => P_HR_NS <= "000000000111" + P_HR_NS396;
				when "01001000010" => P_HR_NS <= "000000001011" + P_HR_NS397;
				when "01001000011" => P_HR_NS <= "000000001011" + P_HR_NS398;
				when "01001000100" => P_HR_NS <= "000000000100" + P_HR_NS399;
				when "01001000101" => P_HR_NS <= "000000000100" + P_HR_NS400;
				when "01001000110" => P_HR_NS <= "000000010010" + P_HR_NS401;
				when "01001000111" => P_HR_NS <= "000000001110" + P_HR_NS402;
				when "01001001000" => P_HR_NS <= "000000011001" + P_HR_NS403;
				when "01001001001" => P_HR_NS <= "000000001110" + P_HR_NS404;
				when "01001001010" => P_HR_NS <= "000000000100" + P_HR_NS405;
				when "01001001011" => P_HR_NS <= "000000000111" + P_HR_NS406;
				when "01001001100" => P_HR_NS <= "000000000100" + P_HR_NS407;
				when "01001001101" => P_HR_NS <= "000000010010" + P_HR_NS408;
				when "01001001111" => P_HR_NS <= "000000000100" + P_HR_NS409;
				when "01001010000" => P_HR_NS <= "000000000100" + P_HR_NS410;
				when "01001010001" => P_HR_NS <= "000000001011" + P_HR_NS411;
				when "01001010010" => P_HR_NS <= "000000001011" + P_HR_NS412;
				when "01001010100" => P_HR_NS <= "000000001011" + P_HR_NS413;
				when "01001010101" => P_HR_NS <= "000000001011" + P_HR_NS414;
				when "01001010110" => P_HR_NS <= "000000000111" + P_HR_NS415;
				when "01001010111" => P_HR_NS <= "000000000100" + P_HR_NS416;
				when "01001011000" => P_HR_NS <= "000000001011" + P_HR_NS417;
				when "01001011001" => P_HR_NS <= "000000001011" + P_HR_NS418;
				when "01001011010" => P_HR_NS <= "000000000100" + P_HR_NS419;
				when "01001011011" => P_HR_NS <= "000000000100" + P_HR_NS420;
				when "01001011101" => P_HR_NS <= "000000000100" + P_HR_NS421;
				when "01001011110" => P_HR_NS <= "000000000100" + P_HR_NS422;
				when "01001100000" => P_HR_NS <= "000000001011" + P_HR_NS423;
				when "01001100010" => P_HR_NS <= "000000000111" + P_HR_NS424;
				when "01001100011" => P_HR_NS <= "000000000100" + P_HR_NS425;
				when "01001100101" => P_HR_NS <= "000000001011" + P_HR_NS426;
				when "01001100110" => P_HR_NS <= "000000001110" + P_HR_NS427;
				when "01001100111" => P_HR_NS <= "000000000100" + P_HR_NS428;
				when "01001101001" => P_HR_NS <= "000000000100" + P_HR_NS429;
				when "01001101010" => P_HR_NS <= "000000000100" + P_HR_NS430;
				when "01001101100" => P_HR_NS <= "000000000100" + P_HR_NS431;
				when "01001101110" => P_HR_NS <= "000000000100" + P_HR_NS432;
				when "01001101111" => P_HR_NS <= "000000000100" + P_HR_NS433;
				when "01001110011" => P_HR_NS <= "000000000100" + P_HR_NS434;
				when "01001111000" => P_HR_NS <= "000000000111" + P_HR_NS435;
				when "01001111011" => P_HR_NS <= "000000000100" + P_HR_NS436;
				when "01010000000" => P_HR_NS <= "000000000100" + P_HR_NS437;
				when "01010000001" => P_HR_NS <= "000000000100" + P_HR_NS438;
				when "01010000100" => P_HR_NS <= "000000000100" + P_HR_NS439;
				when "01010000110" => P_HR_NS <= "000000000100" + P_HR_NS440;
				when "01010001001" => P_HR_NS <= "000000000100" + P_HR_NS441;
				when "01010001010" => P_HR_NS <= "000000000100" + P_HR_NS442;
				when "01010001100" => P_HR_NS <= "000000000100" + P_HR_NS443;
				when "01010011001" => P_HR_NS <= "000000000100" + P_HR_NS444;
				when "01010011100" => P_HR_NS <= "000000000100" + P_HR_NS445;
				when "01010011111" => P_HR_NS <= "000000000100" + P_HR_NS446;
				when "01010100101" => P_HR_NS <= "000000000100" + P_HR_NS447;
				when "01010101000" => P_HR_NS <= "000000000100" + P_HR_NS448;
				when "01010101010" => P_HR_NS <= "000000000100" + P_HR_NS449;
				when "01010111100" => P_HR_NS <= "000000000100" + P_HR_NS450;
				when "01011000010" => P_HR_NS <= "000000000100" + P_HR_NS451;
				when "01011100100" => P_HR_NS <= "000000000100" + P_HR_NS452;
				when "01011101001" => P_HR_NS <= "000000000100" + P_HR_NS453;
				when "10100101011" => P_HR_NS <= "000000000100" + P_HR_NS454;
				when "10101100111" => P_HR_NS <= "000000000100" + P_HR_NS455;
				when others            => P_HR_NS <= "000000000001";
			end case;

			case eda is
				when "0000010" => P_EDA_NS <= "000000000001" + P_EDA_NS1;
				when "0000011" => P_EDA_NS <= "000000000010" + P_EDA_NS2;
				when "0000100" => P_EDA_NS <= "000110100000" + P_EDA_NS3;
				when "0000101" => P_EDA_NS <= "000111101111" + P_EDA_NS4;
				when "0000110" => P_EDA_NS <= "001100010010" + P_EDA_NS5;
				when "0000111" => P_EDA_NS <= "001010010101" + P_EDA_NS6;
				when "0001000" => P_EDA_NS <= "000000111100" + P_EDA_NS7;
				when "0001001" => P_EDA_NS <= "000110010101" + P_EDA_NS8;
				when "0001010" => P_EDA_NS <= "000100100000" + P_EDA_NS9;
				when "0001011" => P_EDA_NS <= "000100001000" + P_EDA_NS10;
				when "0001100" => P_EDA_NS <= "000100001000" + P_EDA_NS11;
				when "0001101" => P_EDA_NS <= "000010101001" + P_EDA_NS12;
				when "0001110" => P_EDA_NS <= "000001110111" + P_EDA_NS13;
				when "0001111" => P_EDA_NS <= "000001011001" + P_EDA_NS14;
				when "0010000" => P_EDA_NS <= "000001001011" + P_EDA_NS15;
				when "0010001" => P_EDA_NS <= "000001000101" + P_EDA_NS16;
				when "0010010" => P_EDA_NS <= "000001000001" + P_EDA_NS17;
				when "0010011" => P_EDA_NS <= "000000110110" + P_EDA_NS18;
				when "0010100" => P_EDA_NS <= "000000101111" + P_EDA_NS19;
				when "0010101" => P_EDA_NS <= "000000101011" + P_EDA_NS20;
				when "0010110" => P_EDA_NS <= "000000100101" + P_EDA_NS21;
				when "0010111" => P_EDA_NS <= "000000100001" + P_EDA_NS22;
				when "0011000" => P_EDA_NS <= "000000011111" + P_EDA_NS23;
				when "0011001" => P_EDA_NS <= "000000011011" + P_EDA_NS24;
				when "0011010" => P_EDA_NS <= "000000011110" + P_EDA_NS25;
				when "0011011" => P_EDA_NS <= "000000110001" + P_EDA_NS26;
				when "0011100" => P_EDA_NS <= "000000011100" + P_EDA_NS27;
				when "0011101" => P_EDA_NS <= "000000011001" + P_EDA_NS28;
				when "0011110" => P_EDA_NS <= "000000011110" + P_EDA_NS29;
				when "0011111" => P_EDA_NS <= "000000011010" + P_EDA_NS30;
				when "0100000" => P_EDA_NS <= "000000011000" + P_EDA_NS31;
				when "0100001" => P_EDA_NS <= "000000010010" + P_EDA_NS32;
				when "0100010" => P_EDA_NS <= "000000010100" + P_EDA_NS33;
				when "0100011" => P_EDA_NS <= "000000010011" + P_EDA_NS34;
				when "0100100" => P_EDA_NS <= "000000010011" + P_EDA_NS35;
				when "0100101" => P_EDA_NS <= "000000010011" + P_EDA_NS36;
				when "0100110" => P_EDA_NS <= "000000011110" + P_EDA_NS37;
				when "0100111" => P_EDA_NS <= "000000001111" + P_EDA_NS38;
				when "0101000" => P_EDA_NS <= "000000001100" + P_EDA_NS39;
				when "0101001" => P_EDA_NS <= "000000011000" + P_EDA_NS40;
				when "0101010" => P_EDA_NS <= "000000001010" + P_EDA_NS41;
				when "0101011" => P_EDA_NS <= "000000001000" + P_EDA_NS42;
				when "0101100" => P_EDA_NS <= "000000000101" + P_EDA_NS43;
				when "0101101" => P_EDA_NS <= "000000000011" + P_EDA_NS44;
				when "0101110" => P_EDA_NS <= "000000000010" + P_EDA_NS45;
				when "0110010" => P_EDA_NS <= "000000000010" + P_EDA_NS46;
				when "0110011" => P_EDA_NS <= "000000000010" + P_EDA_NS47;
				when "0110100" => P_EDA_NS <= "001000100111" + P_EDA_NS48;
				when "0110101" => P_EDA_NS <= "001011101100" + P_EDA_NS49;
				when "0110110" => P_EDA_NS <= "000100101001" + P_EDA_NS50;
				when "0110111" => P_EDA_NS <= "000001011011" + P_EDA_NS51;
				when "0111000" => P_EDA_NS <= "000010100111" + P_EDA_NS52;
				when "0111001" => P_EDA_NS <= "001111010101" + P_EDA_NS53;
				when "0111010" => P_EDA_NS <= "000101010001" + P_EDA_NS54;
				when "0111011" => P_EDA_NS <= "000100101001" + P_EDA_NS55;
				when "0111100" => P_EDA_NS <= "000101000001" + P_EDA_NS56;
				when "0111101" => P_EDA_NS <= "000000111110" + P_EDA_NS57;
				when "0111110" => P_EDA_NS <= "000011000110" + P_EDA_NS58;
				when "0111111" => P_EDA_NS <= "000100000000" + P_EDA_NS59;
				when "1000000" => P_EDA_NS <= "000010111010" + P_EDA_NS60;
				when "1000001" => P_EDA_NS <= "000011100000" + P_EDA_NS61;
				when "1000010" => P_EDA_NS <= "000010110100" + P_EDA_NS62;
				when "1000011" => P_EDA_NS <= "000000010111" + P_EDA_NS63;
				when "1000100" => P_EDA_NS <= "000000100000" + P_EDA_NS64;
				when "1000101" => P_EDA_NS <= "000000100101" + P_EDA_NS65;
				when "1000110" => P_EDA_NS <= "000001001101" + P_EDA_NS66;
				when "1000111" => P_EDA_NS <= "000000010000" + P_EDA_NS67;
				when others    => P_EDA_NS <= "000000000001";
			end case;
			not_stress_score <= P_TEMP_NS * P_NOT_STRESS * P_EDA_NS * P_HR_NS;
			
			--not_stress_score <= P_TEMP_NS * P_NOT_STRESS * P_EDA_NS * P_HR_NS;
		elsif (state = TRAINING_NS) then
			
			case temp is
				when "011100000" => P_TEMP_NS1   <= P_TEMP_NS1 + "111101000";
				when "011100001" => P_TEMP_NS2   <= P_TEMP_NS2 + "111101000";
				when "011100010" => P_TEMP_NS3   <= P_TEMP_NS3 + "111101000";
				when "011100011" => P_TEMP_NS4   <= P_TEMP_NS4 + "111101000";
				when "011100100" => P_TEMP_NS5   <= P_TEMP_NS5 + "111101000";
				when "011100101" => P_TEMP_NS6   <= P_TEMP_NS6 + "111101000";
				when "011100110" => P_TEMP_NS7   <= P_TEMP_NS7 + "111101000";
				when "011100111" => P_TEMP_NS8   <= P_TEMP_NS8 + "111101000";
				when "011101000" => P_TEMP_NS9   <= P_TEMP_NS9 + "111101000";
				when "011101001" => P_TEMP_NS10 <= P_TEMP_NS10 + "111101000";
				when "011101010" => P_TEMP_NS11 <= P_TEMP_NS11 + "111101000";
				when "011101011" => P_TEMP_NS12 <= P_TEMP_NS12 + "111101000";
				when "011101100" => P_TEMP_NS13 <= P_TEMP_NS13 + "111101000";
				when "011101101" => P_TEMP_NS14 <= P_TEMP_NS14 + "111101000";
				when "011101110" => P_TEMP_NS15 <= P_TEMP_NS15 + "111101000";
				when "011101111" => P_TEMP_NS16 <= P_TEMP_NS16 + "111101000";
				when "011110000" => P_TEMP_NS17 <= P_TEMP_NS17 + "111101000";
				when "011110001" => P_TEMP_NS18 <= P_TEMP_NS18 + "111101000";
				when "011110010" => P_TEMP_NS19 <= P_TEMP_NS19 + "111101000";
				when "011110011" => P_TEMP_NS20 <= P_TEMP_NS20 + "111101000";
				when "011110100" => P_TEMP_NS21 <= P_TEMP_NS21 + "111101000";
				when "011110101" => P_TEMP_NS22 <= P_TEMP_NS22 + "111101000";
				when "011110110" => P_TEMP_NS23 <= P_TEMP_NS23 + "111101000";
				when "011110111" => P_TEMP_NS24 <= P_TEMP_NS24 + "111101000";
				when "011111000" => P_TEMP_NS25 <= P_TEMP_NS25 + "111101000";
				when "011111001" => P_TEMP_NS26 <= P_TEMP_NS26 + "111101000";
				when "011111010" => P_TEMP_NS27 <= P_TEMP_NS27 + "111101000";
				when "011111011" => P_TEMP_NS28 <= P_TEMP_NS28 + "111101000";
				when "011111100" => P_TEMP_NS29 <= P_TEMP_NS29 + "111101000";
				when "011111101" => P_TEMP_NS30 <= P_TEMP_NS30 + "111101000";
				when "011111110" => P_TEMP_NS31 <= P_TEMP_NS31 + "111101000";
				when "011111111" => P_TEMP_NS32 <= P_TEMP_NS32 + "111101000";
				when "100000000" => P_TEMP_NS33 <= P_TEMP_NS33 + "111101000";
				when "100000001" => P_TEMP_NS34 <= P_TEMP_NS34 + "111101000";
				when "100000010" => P_TEMP_NS35 <= P_TEMP_NS35 + "111101000";
				when "100000011" => P_TEMP_NS36 <= P_TEMP_NS36 + "111101000";
				when "100000100" => P_TEMP_NS37 <= P_TEMP_NS37 + "111101000";
				when "100000101" => P_TEMP_NS38 <= P_TEMP_NS38 + "111101000";
				when "100000110" => P_TEMP_NS39 <= P_TEMP_NS39 + "111101000";
				when "100000111" => P_TEMP_NS40 <= P_TEMP_NS40 + "111101000";
				when "100001000" => P_TEMP_NS41 <= P_TEMP_NS41 + "111101000";
				when "100001001" => P_TEMP_NS42 <= P_TEMP_NS42 + "111101000";
				when "100001010" => P_TEMP_NS43 <= P_TEMP_NS43 + "111101000";
				when "100001011" => P_TEMP_NS44 <= P_TEMP_NS44 + "111101000";
				when "100001100" => P_TEMP_NS45 <= P_TEMP_NS45 + "111101000";
				when "100001101" => P_TEMP_NS46 <= P_TEMP_NS46 + "111101000";
				when "100001110" => P_TEMP_NS47 <= P_TEMP_NS47 + "111101000";
				when "100001111" => P_TEMP_NS48 <= P_TEMP_NS48 + "111101000";
				when "100010000" => P_TEMP_NS49 <= P_TEMP_NS49 + "111101000";
				when "100010001" => P_TEMP_NS50 <= P_TEMP_NS50 + "111101000";
				when "100010010" => P_TEMP_NS51 <= P_TEMP_NS51 + "111101000";
				when "100010011" => P_TEMP_NS52 <= P_TEMP_NS52 + "111101000";
				when  others     => null;
			end case;	

			
		else -- in training mode
			not_stress_score <= (others => '0');
			P_TEMP_NS <= (others => '0'); 
			P_EDA_NS <= (others => '0');
			P_HR_NS <= (others => '0');
		end if;
	   end if;
	end process;
	


end behavioral;